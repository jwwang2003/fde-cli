
module top ( clk, clk_30M, rst, nReset, i_wr, i_wdata, i_rd, o_rdata, o_rempty, 
        o_wfull, fifo_1_w_full );
  input [7:0] i_wdata;
  output [7:0] o_rdata;
  input clk, clk_30M, rst, nReset, i_wr, i_rd;
  output o_rempty, o_wfull, fifo_1_w_full;
  wire   active, rd_fifo_empty, N2, \fifo_write/rempty_next ,
         \fifo_write/rgraynext[0] , \fifo_write/rgraynext[1] ,
         \fifo_write/rgraynext[2] , \fifo_write/rgraynext[3] ,
         \fifo_write/rgraynext[4] , \fifo_write/rbinnext[0] ,
         \fifo_write/rbinnext[1] , \fifo_write/rbinnext[2] ,
         \fifo_write/rbinnext[3] , \fifo_write/rbinnext[4] ,
         \fifo_write/rbinnext[5] , \fifo_write/rbin[0] , \fifo_write/rbin[1] ,
         \fifo_write/rbin[2] , \fifo_write/rbin[3] , \fifo_write/rbin[4] ,
         \fifo_write/mem[0][7] , \fifo_write/mem[0][6] ,
         \fifo_write/mem[0][5] , \fifo_write/mem[0][4] ,
         \fifo_write/mem[0][3] , \fifo_write/mem[0][2] ,
         \fifo_write/mem[0][1] , \fifo_write/mem[0][0] ,
         \fifo_write/mem[1][7] , \fifo_write/mem[1][6] ,
         \fifo_write/mem[1][5] , \fifo_write/mem[1][4] ,
         \fifo_write/mem[1][3] , \fifo_write/mem[1][2] ,
         \fifo_write/mem[1][1] , \fifo_write/mem[1][0] ,
         \fifo_write/mem[2][7] , \fifo_write/mem[2][6] ,
         \fifo_write/mem[2][5] , \fifo_write/mem[2][4] ,
         \fifo_write/mem[2][3] , \fifo_write/mem[2][2] ,
         \fifo_write/mem[2][1] , \fifo_write/mem[2][0] ,
         \fifo_write/mem[3][7] , \fifo_write/mem[3][6] ,
         \fifo_write/mem[3][5] , \fifo_write/mem[3][4] ,
         \fifo_write/mem[3][3] , \fifo_write/mem[3][2] ,
         \fifo_write/mem[3][1] , \fifo_write/mem[3][0] ,
         \fifo_write/mem[4][7] , \fifo_write/mem[4][6] ,
         \fifo_write/mem[4][5] , \fifo_write/mem[4][4] ,
         \fifo_write/mem[4][3] , \fifo_write/mem[4][2] ,
         \fifo_write/mem[4][1] , \fifo_write/mem[4][0] ,
         \fifo_write/mem[5][7] , \fifo_write/mem[5][6] ,
         \fifo_write/mem[5][5] , \fifo_write/mem[5][4] ,
         \fifo_write/mem[5][3] , \fifo_write/mem[5][2] ,
         \fifo_write/mem[5][1] , \fifo_write/mem[5][0] ,
         \fifo_write/mem[6][7] , \fifo_write/mem[6][6] ,
         \fifo_write/mem[6][5] , \fifo_write/mem[6][4] ,
         \fifo_write/mem[6][3] , \fifo_write/mem[6][2] ,
         \fifo_write/mem[6][1] , \fifo_write/mem[6][0] ,
         \fifo_write/mem[7][7] , \fifo_write/mem[7][6] ,
         \fifo_write/mem[7][5] , \fifo_write/mem[7][4] ,
         \fifo_write/mem[7][3] , \fifo_write/mem[7][2] ,
         \fifo_write/mem[7][1] , \fifo_write/mem[7][0] ,
         \fifo_write/mem[8][7] , \fifo_write/mem[8][6] ,
         \fifo_write/mem[8][5] , \fifo_write/mem[8][4] ,
         \fifo_write/mem[8][3] , \fifo_write/mem[8][2] ,
         \fifo_write/mem[8][1] , \fifo_write/mem[8][0] ,
         \fifo_write/mem[9][7] , \fifo_write/mem[9][6] ,
         \fifo_write/mem[9][5] , \fifo_write/mem[9][4] ,
         \fifo_write/mem[9][3] , \fifo_write/mem[9][2] ,
         \fifo_write/mem[9][1] , \fifo_write/mem[9][0] ,
         \fifo_write/mem[10][7] , \fifo_write/mem[10][6] ,
         \fifo_write/mem[10][5] , \fifo_write/mem[10][4] ,
         \fifo_write/mem[10][3] , \fifo_write/mem[10][2] ,
         \fifo_write/mem[10][1] , \fifo_write/mem[10][0] ,
         \fifo_write/mem[11][7] , \fifo_write/mem[11][6] ,
         \fifo_write/mem[11][5] , \fifo_write/mem[11][4] ,
         \fifo_write/mem[11][3] , \fifo_write/mem[11][2] ,
         \fifo_write/mem[11][1] , \fifo_write/mem[11][0] ,
         \fifo_write/mem[12][7] , \fifo_write/mem[12][6] ,
         \fifo_write/mem[12][5] , \fifo_write/mem[12][4] ,
         \fifo_write/mem[12][3] , \fifo_write/mem[12][2] ,
         \fifo_write/mem[12][1] , \fifo_write/mem[12][0] ,
         \fifo_write/mem[13][7] , \fifo_write/mem[13][6] ,
         \fifo_write/mem[13][5] , \fifo_write/mem[13][4] ,
         \fifo_write/mem[13][3] , \fifo_write/mem[13][2] ,
         \fifo_write/mem[13][1] , \fifo_write/mem[13][0] ,
         \fifo_write/mem[14][7] , \fifo_write/mem[14][6] ,
         \fifo_write/mem[14][5] , \fifo_write/mem[14][4] ,
         \fifo_write/mem[14][3] , \fifo_write/mem[14][2] ,
         \fifo_write/mem[14][1] , \fifo_write/mem[14][0] ,
         \fifo_write/mem[15][7] , \fifo_write/mem[15][6] ,
         \fifo_write/mem[15][5] , \fifo_write/mem[15][4] ,
         \fifo_write/mem[15][3] , \fifo_write/mem[15][2] ,
         \fifo_write/mem[15][1] , \fifo_write/mem[15][0] ,
         \fifo_write/mem[16][7] , \fifo_write/mem[16][6] ,
         \fifo_write/mem[16][5] , \fifo_write/mem[16][4] ,
         \fifo_write/mem[16][3] , \fifo_write/mem[16][2] ,
         \fifo_write/mem[16][1] , \fifo_write/mem[16][0] ,
         \fifo_write/mem[17][7] , \fifo_write/mem[17][6] ,
         \fifo_write/mem[17][5] , \fifo_write/mem[17][4] ,
         \fifo_write/mem[17][3] , \fifo_write/mem[17][2] ,
         \fifo_write/mem[17][1] , \fifo_write/mem[17][0] ,
         \fifo_write/mem[18][7] , \fifo_write/mem[18][6] ,
         \fifo_write/mem[18][5] , \fifo_write/mem[18][4] ,
         \fifo_write/mem[18][3] , \fifo_write/mem[18][2] ,
         \fifo_write/mem[18][1] , \fifo_write/mem[18][0] ,
         \fifo_write/mem[19][7] , \fifo_write/mem[19][6] ,
         \fifo_write/mem[19][5] , \fifo_write/mem[19][4] ,
         \fifo_write/mem[19][3] , \fifo_write/mem[19][2] ,
         \fifo_write/mem[19][1] , \fifo_write/mem[19][0] ,
         \fifo_write/mem[20][7] , \fifo_write/mem[20][6] ,
         \fifo_write/mem[20][5] , \fifo_write/mem[20][4] ,
         \fifo_write/mem[20][3] , \fifo_write/mem[20][2] ,
         \fifo_write/mem[20][1] , \fifo_write/mem[20][0] ,
         \fifo_write/mem[21][7] , \fifo_write/mem[21][6] ,
         \fifo_write/mem[21][5] , \fifo_write/mem[21][4] ,
         \fifo_write/mem[21][3] , \fifo_write/mem[21][2] ,
         \fifo_write/mem[21][1] , \fifo_write/mem[21][0] ,
         \fifo_write/mem[22][7] , \fifo_write/mem[22][6] ,
         \fifo_write/mem[22][5] , \fifo_write/mem[22][4] ,
         \fifo_write/mem[22][3] , \fifo_write/mem[22][2] ,
         \fifo_write/mem[22][1] , \fifo_write/mem[22][0] ,
         \fifo_write/mem[23][7] , \fifo_write/mem[23][6] ,
         \fifo_write/mem[23][5] , \fifo_write/mem[23][4] ,
         \fifo_write/mem[23][3] , \fifo_write/mem[23][2] ,
         \fifo_write/mem[23][1] , \fifo_write/mem[23][0] ,
         \fifo_write/mem[24][7] , \fifo_write/mem[24][6] ,
         \fifo_write/mem[24][5] , \fifo_write/mem[24][4] ,
         \fifo_write/mem[24][3] , \fifo_write/mem[24][2] ,
         \fifo_write/mem[24][1] , \fifo_write/mem[24][0] ,
         \fifo_write/mem[25][7] , \fifo_write/mem[25][6] ,
         \fifo_write/mem[25][5] , \fifo_write/mem[25][4] ,
         \fifo_write/mem[25][3] , \fifo_write/mem[25][2] ,
         \fifo_write/mem[25][1] , \fifo_write/mem[25][0] ,
         \fifo_write/mem[26][7] , \fifo_write/mem[26][6] ,
         \fifo_write/mem[26][5] , \fifo_write/mem[26][4] ,
         \fifo_write/mem[26][3] , \fifo_write/mem[26][2] ,
         \fifo_write/mem[26][1] , \fifo_write/mem[26][0] ,
         \fifo_write/mem[27][7] , \fifo_write/mem[27][6] ,
         \fifo_write/mem[27][5] , \fifo_write/mem[27][4] ,
         \fifo_write/mem[27][3] , \fifo_write/mem[27][2] ,
         \fifo_write/mem[27][1] , \fifo_write/mem[27][0] ,
         \fifo_write/mem[28][7] , \fifo_write/mem[28][6] ,
         \fifo_write/mem[28][5] , \fifo_write/mem[28][4] ,
         \fifo_write/mem[28][3] , \fifo_write/mem[28][2] ,
         \fifo_write/mem[28][1] , \fifo_write/mem[28][0] ,
         \fifo_write/mem[29][7] , \fifo_write/mem[29][6] ,
         \fifo_write/mem[29][5] , \fifo_write/mem[29][4] ,
         \fifo_write/mem[29][3] , \fifo_write/mem[29][2] ,
         \fifo_write/mem[29][1] , \fifo_write/mem[29][0] ,
         \fifo_write/mem[30][7] , \fifo_write/mem[30][6] ,
         \fifo_write/mem[30][5] , \fifo_write/mem[30][4] ,
         \fifo_write/mem[30][3] , \fifo_write/mem[30][2] ,
         \fifo_write/mem[30][1] , \fifo_write/mem[30][0] ,
         \fifo_write/mem[31][7] , \fifo_write/mem[31][6] ,
         \fifo_write/mem[31][5] , \fifo_write/mem[31][4] ,
         \fifo_write/mem[31][3] , \fifo_write/mem[31][2] ,
         \fifo_write/mem[31][1] , \fifo_write/mem[31][0] ,
         \fifo_write/wfull_next , \fifo_write/waddr[0] , \fifo_write/waddr[1] ,
         \fifo_write/waddr[2] , \fifo_write/waddr[3] , \fifo_write/waddr[4] ,
         \fifo_write/wgraynext[0] , \fifo_write/wgraynext[1] ,
         \fifo_write/wgraynext[2] , \fifo_write/wgraynext[3] ,
         \fifo_write/wgraynext[4] , \fifo_write/wbinnext[0] ,
         \fifo_write/wbinnext[1] , \fifo_write/wbinnext[2] ,
         \fifo_write/wbinnext[3] , \fifo_write/wbinnext[4] ,
         \fifo_write/wbinnext[5] , \fifo_read/rempty_next ,
         \fifo_read/rgraynext[0] , \fifo_read/rgraynext[1] ,
         \fifo_read/rgraynext[2] , \fifo_read/rgraynext[3] ,
         \fifo_read/rgraynext[4] , \fifo_read/rbinnext[0] ,
         \fifo_read/rbinnext[1] , \fifo_read/rbinnext[2] ,
         \fifo_read/rbinnext[3] , \fifo_read/rbinnext[4] ,
         \fifo_read/rbinnext[5] , \fifo_read/rbin[0] , \fifo_read/rbin[1] ,
         \fifo_read/rbin[2] , \fifo_read/rbin[3] , \fifo_read/rbin[4] ,
         \fifo_read/mem[0][7] , \fifo_read/mem[0][6] , \fifo_read/mem[0][5] ,
         \fifo_read/mem[0][4] , \fifo_read/mem[0][3] , \fifo_read/mem[0][2] ,
         \fifo_read/mem[0][1] , \fifo_read/mem[0][0] , \fifo_read/mem[1][7] ,
         \fifo_read/mem[1][6] , \fifo_read/mem[1][5] , \fifo_read/mem[1][4] ,
         \fifo_read/mem[1][3] , \fifo_read/mem[1][2] , \fifo_read/mem[1][1] ,
         \fifo_read/mem[1][0] , \fifo_read/mem[2][7] , \fifo_read/mem[2][6] ,
         \fifo_read/mem[2][5] , \fifo_read/mem[2][4] , \fifo_read/mem[2][3] ,
         \fifo_read/mem[2][2] , \fifo_read/mem[2][1] , \fifo_read/mem[2][0] ,
         \fifo_read/mem[3][7] , \fifo_read/mem[3][6] , \fifo_read/mem[3][5] ,
         \fifo_read/mem[3][4] , \fifo_read/mem[3][3] , \fifo_read/mem[3][2] ,
         \fifo_read/mem[3][1] , \fifo_read/mem[3][0] , \fifo_read/mem[4][7] ,
         \fifo_read/mem[4][6] , \fifo_read/mem[4][5] , \fifo_read/mem[4][4] ,
         \fifo_read/mem[4][3] , \fifo_read/mem[4][2] , \fifo_read/mem[4][1] ,
         \fifo_read/mem[4][0] , \fifo_read/mem[5][7] , \fifo_read/mem[5][6] ,
         \fifo_read/mem[5][5] , \fifo_read/mem[5][4] , \fifo_read/mem[5][3] ,
         \fifo_read/mem[5][2] , \fifo_read/mem[5][1] , \fifo_read/mem[5][0] ,
         \fifo_read/mem[6][7] , \fifo_read/mem[6][6] , \fifo_read/mem[6][5] ,
         \fifo_read/mem[6][4] , \fifo_read/mem[6][3] , \fifo_read/mem[6][2] ,
         \fifo_read/mem[6][1] , \fifo_read/mem[6][0] , \fifo_read/mem[7][7] ,
         \fifo_read/mem[7][6] , \fifo_read/mem[7][5] , \fifo_read/mem[7][4] ,
         \fifo_read/mem[7][3] , \fifo_read/mem[7][2] , \fifo_read/mem[7][1] ,
         \fifo_read/mem[7][0] , \fifo_read/mem[8][7] , \fifo_read/mem[8][6] ,
         \fifo_read/mem[8][5] , \fifo_read/mem[8][4] , \fifo_read/mem[8][3] ,
         \fifo_read/mem[8][2] , \fifo_read/mem[8][1] , \fifo_read/mem[8][0] ,
         \fifo_read/mem[9][7] , \fifo_read/mem[9][6] , \fifo_read/mem[9][5] ,
         \fifo_read/mem[9][4] , \fifo_read/mem[9][3] , \fifo_read/mem[9][2] ,
         \fifo_read/mem[9][1] , \fifo_read/mem[9][0] , \fifo_read/mem[10][7] ,
         \fifo_read/mem[10][6] , \fifo_read/mem[10][5] ,
         \fifo_read/mem[10][4] , \fifo_read/mem[10][3] ,
         \fifo_read/mem[10][2] , \fifo_read/mem[10][1] ,
         \fifo_read/mem[10][0] , \fifo_read/mem[11][7] ,
         \fifo_read/mem[11][6] , \fifo_read/mem[11][5] ,
         \fifo_read/mem[11][4] , \fifo_read/mem[11][3] ,
         \fifo_read/mem[11][2] , \fifo_read/mem[11][1] ,
         \fifo_read/mem[11][0] , \fifo_read/mem[12][7] ,
         \fifo_read/mem[12][6] , \fifo_read/mem[12][5] ,
         \fifo_read/mem[12][4] , \fifo_read/mem[12][3] ,
         \fifo_read/mem[12][2] , \fifo_read/mem[12][1] ,
         \fifo_read/mem[12][0] , \fifo_read/mem[13][7] ,
         \fifo_read/mem[13][6] , \fifo_read/mem[13][5] ,
         \fifo_read/mem[13][4] , \fifo_read/mem[13][3] ,
         \fifo_read/mem[13][2] , \fifo_read/mem[13][1] ,
         \fifo_read/mem[13][0] , \fifo_read/mem[14][7] ,
         \fifo_read/mem[14][6] , \fifo_read/mem[14][5] ,
         \fifo_read/mem[14][4] , \fifo_read/mem[14][3] ,
         \fifo_read/mem[14][2] , \fifo_read/mem[14][1] ,
         \fifo_read/mem[14][0] , \fifo_read/mem[15][7] ,
         \fifo_read/mem[15][6] , \fifo_read/mem[15][5] ,
         \fifo_read/mem[15][4] , \fifo_read/mem[15][3] ,
         \fifo_read/mem[15][2] , \fifo_read/mem[15][1] ,
         \fifo_read/mem[15][0] , \fifo_read/mem[16][7] ,
         \fifo_read/mem[16][6] , \fifo_read/mem[16][5] ,
         \fifo_read/mem[16][4] , \fifo_read/mem[16][3] ,
         \fifo_read/mem[16][2] , \fifo_read/mem[16][1] ,
         \fifo_read/mem[16][0] , \fifo_read/mem[17][7] ,
         \fifo_read/mem[17][6] , \fifo_read/mem[17][5] ,
         \fifo_read/mem[17][4] , \fifo_read/mem[17][3] ,
         \fifo_read/mem[17][2] , \fifo_read/mem[17][1] ,
         \fifo_read/mem[17][0] , \fifo_read/mem[18][7] ,
         \fifo_read/mem[18][6] , \fifo_read/mem[18][5] ,
         \fifo_read/mem[18][4] , \fifo_read/mem[18][3] ,
         \fifo_read/mem[18][2] , \fifo_read/mem[18][1] ,
         \fifo_read/mem[18][0] , \fifo_read/mem[19][7] ,
         \fifo_read/mem[19][6] , \fifo_read/mem[19][5] ,
         \fifo_read/mem[19][4] , \fifo_read/mem[19][3] ,
         \fifo_read/mem[19][2] , \fifo_read/mem[19][1] ,
         \fifo_read/mem[19][0] , \fifo_read/mem[20][7] ,
         \fifo_read/mem[20][6] , \fifo_read/mem[20][5] ,
         \fifo_read/mem[20][4] , \fifo_read/mem[20][3] ,
         \fifo_read/mem[20][2] , \fifo_read/mem[20][1] ,
         \fifo_read/mem[20][0] , \fifo_read/mem[21][7] ,
         \fifo_read/mem[21][6] , \fifo_read/mem[21][5] ,
         \fifo_read/mem[21][4] , \fifo_read/mem[21][3] ,
         \fifo_read/mem[21][2] , \fifo_read/mem[21][1] ,
         \fifo_read/mem[21][0] , \fifo_read/mem[22][7] ,
         \fifo_read/mem[22][6] , \fifo_read/mem[22][5] ,
         \fifo_read/mem[22][4] , \fifo_read/mem[22][3] ,
         \fifo_read/mem[22][2] , \fifo_read/mem[22][1] ,
         \fifo_read/mem[22][0] , \fifo_read/mem[23][7] ,
         \fifo_read/mem[23][6] , \fifo_read/mem[23][5] ,
         \fifo_read/mem[23][4] , \fifo_read/mem[23][3] ,
         \fifo_read/mem[23][2] , \fifo_read/mem[23][1] ,
         \fifo_read/mem[23][0] , \fifo_read/mem[24][7] ,
         \fifo_read/mem[24][6] , \fifo_read/mem[24][5] ,
         \fifo_read/mem[24][4] , \fifo_read/mem[24][3] ,
         \fifo_read/mem[24][2] , \fifo_read/mem[24][1] ,
         \fifo_read/mem[24][0] , \fifo_read/mem[25][7] ,
         \fifo_read/mem[25][6] , \fifo_read/mem[25][5] ,
         \fifo_read/mem[25][4] , \fifo_read/mem[25][3] ,
         \fifo_read/mem[25][2] , \fifo_read/mem[25][1] ,
         \fifo_read/mem[25][0] , \fifo_read/mem[26][7] ,
         \fifo_read/mem[26][6] , \fifo_read/mem[26][5] ,
         \fifo_read/mem[26][4] , \fifo_read/mem[26][3] ,
         \fifo_read/mem[26][2] , \fifo_read/mem[26][1] ,
         \fifo_read/mem[26][0] , \fifo_read/mem[27][7] ,
         \fifo_read/mem[27][6] , \fifo_read/mem[27][5] ,
         \fifo_read/mem[27][4] , \fifo_read/mem[27][3] ,
         \fifo_read/mem[27][2] , \fifo_read/mem[27][1] ,
         \fifo_read/mem[27][0] , \fifo_read/mem[28][7] ,
         \fifo_read/mem[28][6] , \fifo_read/mem[28][5] ,
         \fifo_read/mem[28][4] , \fifo_read/mem[28][3] ,
         \fifo_read/mem[28][2] , \fifo_read/mem[28][1] ,
         \fifo_read/mem[28][0] , \fifo_read/mem[29][7] ,
         \fifo_read/mem[29][6] , \fifo_read/mem[29][5] ,
         \fifo_read/mem[29][4] , \fifo_read/mem[29][3] ,
         \fifo_read/mem[29][2] , \fifo_read/mem[29][1] ,
         \fifo_read/mem[29][0] , \fifo_read/mem[30][7] ,
         \fifo_read/mem[30][6] , \fifo_read/mem[30][5] ,
         \fifo_read/mem[30][4] , \fifo_read/mem[30][3] ,
         \fifo_read/mem[30][2] , \fifo_read/mem[30][1] ,
         \fifo_read/mem[30][0] , \fifo_read/mem[31][7] ,
         \fifo_read/mem[31][6] , \fifo_read/mem[31][5] ,
         \fifo_read/mem[31][4] , \fifo_read/mem[31][3] ,
         \fifo_read/mem[31][2] , \fifo_read/mem[31][1] ,
         \fifo_read/mem[31][0] , \fifo_read/wfull_next , \fifo_read/waddr[0] ,
         \fifo_read/waddr[1] , \fifo_read/waddr[2] , \fifo_read/waddr[3] ,
         \fifo_read/waddr[4] , \fifo_read/wgraynext[0] ,
         \fifo_read/wgraynext[1] , \fifo_read/wgraynext[2] ,
         \fifo_read/wgraynext[3] , \fifo_read/wgraynext[4] ,
         \fifo_read/wbinnext[0] , \fifo_read/wbinnext[1] ,
         \fifo_read/wbinnext[2] , \fifo_read/wbinnext[3] ,
         \fifo_read/wbinnext[4] , \fifo_read/wbinnext[5] , n185, n186, n187,
         n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198,
         n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209,
         n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220,
         n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231,
         n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242,
         n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253,
         n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, n264,
         n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, n275,
         n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286,
         n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297,
         n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308,
         n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319,
         n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330,
         n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341,
         n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352,
         n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
         n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374,
         n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385,
         n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396,
         n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407,
         n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418,
         n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429,
         n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440,
         n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451,
         n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462,
         n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473,
         n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484,
         n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495,
         n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506,
         n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517,
         n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528,
         n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
         n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550,
         n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
         n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572,
         n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583,
         n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594,
         n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605,
         n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616,
         n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627,
         n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638,
         n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649,
         n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660,
         n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671,
         n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682,
         n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693,
         n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704,
         n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715,
         n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726,
         n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737,
         n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748,
         n749, n750, n751, n752, n753, n754, n755, n756, n757, n758, n759,
         n760, n761, n762, n763, n764, n765, n766, n767, n768, n769, n770,
         n771, n772, n773, n774, n775, n776, n777, n778, n779, n780, n781,
         n782, n783, n784, n785, n786, n787, n788, n789, n790, n791, n792,
         n793, n794, n795, n796, n797, n798, n799, n800, n801, n802, n803,
         n804, n805, n806, n807, n808, n809, n810, n811, n812, n813, n814,
         n815, n816, n817, n818, n819, n820, n821, n822, n823, n824, n825,
         n826, n827, n828, n829, n830, n831, n832, n833, n834, n835, n836,
         n837, n838, n839, n840, n841, n842, n843, n844, n845, n846, n847,
         n848, n849, n850, n851, n852, n853, n854, n855, n856, n857, n858,
         n859, n860, n861, n862, n863, n864, n865, n866, n867, n868, n869,
         n870, n871, n872, n873, n874, n875, n876, n877, n878, n879, n880,
         n881, n882, n883, n884, n885, n886, n887, n888, n889, n890, n891,
         n892, n893, n894, n895, n896, n897, n898, n899, n900, n901, n902,
         n903, n904, n905, n906, n907, n908, n909, n910, n911, n912, n913,
         n914, n915, n916, n917, n918, n919, n920, n921, n922, n923, n924,
         n925, n926, n927, n928, n929, n930, n931, n932, n933, n934, n935,
         n936, n937, n938, n939, n940, n941, n942, n943, n944, n945, n946,
         n947, n948, n949, n950, n951, n952, n953, n954, n955, n956, n957,
         n958, n959, n960, n961, n962, n963, n964, n965, n966, n967, n968,
         n969, n970, n971, n972, n973, n974, n975, n976, n977, n978, n979,
         n980, n981, n982, n983, n984, n985, n986, n987, n988, n989, n990,
         n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001,
         n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011,
         n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021,
         n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031,
         n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041,
         n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051,
         n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061,
         n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071,
         n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081,
         n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091,
         n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101,
         n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111,
         n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121,
         n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131,
         n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141,
         n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151,
         n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161,
         n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171,
         n1172, n1173, n1174, n1175, n1176, n1181, n1182, n1183, n1184, n1185,
         n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195,
         n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205,
         n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215,
         n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225,
         n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235,
         n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245,
         n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255,
         n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265,
         n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275,
         n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285,
         n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295,
         n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305,
         n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315,
         n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325,
         n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335,
         n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345,
         n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355,
         n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365,
         n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375,
         n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385,
         n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395,
         n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405,
         n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415,
         n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424, n1425,
         n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434, n1435,
         n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444, n1445,
         n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454, n1455,
         n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464, n1465,
         n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474, n1475,
         n1476, n1477, n1478, n1479, n1480, n1481, n1482, n1483, n1484, n1485,
         n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494, n1495,
         n1496, n1497, n1498, n1499, n1500, n1501, n1502, n1503, n1504, n1505,
         n1506, n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1514, n1515,
         n1516, n1517, n1518;
  wire   [7:0] wdata_to_fifo;
  wire   [5:0] \fifo_write/rq2_wgray ;
  wire   [5:0] \fifo_write/rq1_wgray ;
  wire   [5:0] \fifo_write/wgray ;
  wire   [5:0] \fifo_write/wq2_rgray ;
  wire   [5:0] \fifo_write/rgray ;
  wire   [5:0] \fifo_write/wq1_rgray ;
  wire   [5:0] \fifo_read/rq2_wgray ;
  wire   [5:0] \fifo_read/rq1_wgray ;
  wire   [5:0] \fifo_read/wgray ;
  wire   [5:0] \fifo_read/wq2_rgray ;
  wire   [5:0] \fifo_read/rgray ;
  wire   [5:0] \fifo_read/wq1_rgray ;

  DFFRHQ \fifo_write/wq1_rgray_reg[5]  ( .D(\fifo_write/rgray [5]), .CK(clk), 
        .RN(nReset), .Q(\fifo_write/wq1_rgray [5]) );
  DFFRHQ \fifo_write/wq2_rgray_reg[5]  ( .D(\fifo_write/wq1_rgray [5]), .CK(
        clk), .RN(nReset), .Q(\fifo_write/wq2_rgray [5]) );
  DFFRHQ \fifo_write/o_wfull_reg  ( .D(\fifo_write/wfull_next ), .CK(clk), 
        .RN(nReset), .Q(fifo_1_w_full) );
  DFFRHQ \fifo_write/wbin_reg[0]  ( .D(\fifo_write/wbinnext[0] ), .CK(clk), 
        .RN(nReset), .Q(\fifo_write/waddr[0] ) );
  DFFRHQ \fifo_write/wbin_reg[1]  ( .D(\fifo_write/wbinnext[1] ), .CK(clk), 
        .RN(nReset), .Q(\fifo_write/waddr[1] ) );
  DFFRHQ \fifo_write/wgray_reg[0]  ( .D(\fifo_write/wgraynext[0] ), .CK(clk), 
        .RN(nReset), .Q(\fifo_write/wgray [0]) );
  DFFRHQ \fifo_write/rq1_wgray_reg[0]  ( .D(\fifo_write/wgray [0]), .CK(
        clk_30M), .RN(nReset), .Q(\fifo_write/rq1_wgray [0]) );
  DFFRHQ \fifo_write/rq2_wgray_reg[0]  ( .D(\fifo_write/rq1_wgray [0]), .CK(
        clk_30M), .RN(nReset), .Q(\fifo_write/rq2_wgray [0]) );
  DFFRHQ \fifo_write/wbin_reg[2]  ( .D(\fifo_write/wbinnext[2] ), .CK(clk), 
        .RN(nReset), .Q(\fifo_write/waddr[2] ) );
  DFFRHQ \fifo_write/wgray_reg[1]  ( .D(\fifo_write/wgraynext[1] ), .CK(clk), 
        .RN(nReset), .Q(\fifo_write/wgray [1]) );
  DFFRHQ \fifo_write/rq1_wgray_reg[1]  ( .D(\fifo_write/wgray [1]), .CK(
        clk_30M), .RN(nReset), .Q(\fifo_write/rq1_wgray [1]) );
  DFFRHQ \fifo_write/rq2_wgray_reg[1]  ( .D(\fifo_write/rq1_wgray [1]), .CK(
        clk_30M), .RN(nReset), .Q(\fifo_write/rq2_wgray [1]) );
  DFFRHQ \fifo_write/wbin_reg[3]  ( .D(\fifo_write/wbinnext[3] ), .CK(clk), 
        .RN(nReset), .Q(\fifo_write/waddr[3] ) );
  DFFRHQ \fifo_write/wgray_reg[2]  ( .D(\fifo_write/wgraynext[2] ), .CK(clk), 
        .RN(nReset), .Q(\fifo_write/wgray [2]) );
  DFFRHQ \fifo_write/rq1_wgray_reg[2]  ( .D(\fifo_write/wgray [2]), .CK(
        clk_30M), .RN(nReset), .Q(\fifo_write/rq1_wgray [2]) );
  DFFRHQ \fifo_write/rq2_wgray_reg[2]  ( .D(\fifo_write/rq1_wgray [2]), .CK(
        clk_30M), .RN(nReset), .Q(\fifo_write/rq2_wgray [2]) );
  DFFRHQ \fifo_write/wbin_reg[4]  ( .D(\fifo_write/wbinnext[4] ), .CK(clk), 
        .RN(nReset), .Q(\fifo_write/waddr[4] ) );
  DFFRHQ \fifo_write/wgray_reg[3]  ( .D(\fifo_write/wgraynext[3] ), .CK(clk), 
        .RN(nReset), .Q(\fifo_write/wgray [3]) );
  DFFRHQ \fifo_write/rq1_wgray_reg[3]  ( .D(\fifo_write/wgray [3]), .CK(
        clk_30M), .RN(nReset), .Q(\fifo_write/rq1_wgray [3]) );
  DFFRHQ \fifo_write/rq2_wgray_reg[3]  ( .D(\fifo_write/rq1_wgray [3]), .CK(
        clk_30M), .RN(nReset), .Q(\fifo_write/rq2_wgray [3]) );
  DFFRHQ \fifo_write/wgray_reg[5]  ( .D(\fifo_write/wbinnext[5] ), .CK(clk), 
        .RN(nReset), .Q(\fifo_write/wgray [5]) );
  DFFRHQ \fifo_write/rq1_wgray_reg[5]  ( .D(\fifo_write/wgray [5]), .CK(
        clk_30M), .RN(nReset), .Q(\fifo_write/rq1_wgray [5]) );
  DFFRHQ \fifo_write/rq2_wgray_reg[5]  ( .D(\fifo_write/rq1_wgray [5]), .CK(
        clk_30M), .RN(nReset), .Q(\fifo_write/rq2_wgray [5]) );
  DFFRHQ \fifo_write/wgray_reg[4]  ( .D(\fifo_write/wgraynext[4] ), .CK(clk), 
        .RN(nReset), .Q(\fifo_write/wgray [4]) );
  DFFRHQ \fifo_write/rq1_wgray_reg[4]  ( .D(\fifo_write/wgray [4]), .CK(
        clk_30M), .RN(nReset), .Q(\fifo_write/rq1_wgray [4]) );
  DFFRHQ \fifo_write/rq2_wgray_reg[4]  ( .D(\fifo_write/rq1_wgray [4]), .CK(
        clk_30M), .RN(nReset), .Q(\fifo_write/rq2_wgray [4]) );
  DFFSHQ \fifo_write/o_rempty_reg  ( .D(\fifo_write/rempty_next ), .CK(clk_30M), .SN(nReset), .Q(rd_fifo_empty) );
  DFFRHQ active_reg ( .D(N2), .CK(clk_30M), .RN(nReset), .Q(active) );
  DFFRHQ \fifo_write/rbin_reg[0]  ( .D(\fifo_write/rbinnext[0] ), .CK(clk_30M), 
        .RN(nReset), .Q(\fifo_write/rbin[0] ) );
  DFFRHQ \fifo_write/rbin_reg[1]  ( .D(\fifo_write/rbinnext[1] ), .CK(clk_30M), 
        .RN(nReset), .Q(\fifo_write/rbin[1] ) );
  DFFRHQ \fifo_write/rgray_reg[0]  ( .D(\fifo_write/rgraynext[0] ), .CK(
        clk_30M), .RN(nReset), .Q(\fifo_write/rgray [0]) );
  DFFRHQ \fifo_write/wq1_rgray_reg[0]  ( .D(\fifo_write/rgray [0]), .CK(clk), 
        .RN(nReset), .Q(\fifo_write/wq1_rgray [0]) );
  DFFRHQ \fifo_write/wq2_rgray_reg[0]  ( .D(\fifo_write/wq1_rgray [0]), .CK(
        clk), .RN(nReset), .Q(\fifo_write/wq2_rgray [0]) );
  DFFRHQ \fifo_write/rbin_reg[2]  ( .D(\fifo_write/rbinnext[2] ), .CK(clk_30M), 
        .RN(nReset), .Q(\fifo_write/rbin[2] ) );
  DFFRHQ \fifo_write/rgray_reg[1]  ( .D(\fifo_write/rgraynext[1] ), .CK(
        clk_30M), .RN(nReset), .Q(\fifo_write/rgray [1]) );
  DFFRHQ \fifo_write/wq1_rgray_reg[1]  ( .D(\fifo_write/rgray [1]), .CK(clk), 
        .RN(nReset), .Q(\fifo_write/wq1_rgray [1]) );
  DFFRHQ \fifo_write/wq2_rgray_reg[1]  ( .D(\fifo_write/wq1_rgray [1]), .CK(
        clk), .RN(nReset), .Q(\fifo_write/wq2_rgray [1]) );
  DFFRHQ \fifo_write/rbin_reg[3]  ( .D(\fifo_write/rbinnext[3] ), .CK(clk_30M), 
        .RN(nReset), .Q(\fifo_write/rbin[3] ) );
  DFFRHQ \fifo_write/rgray_reg[2]  ( .D(\fifo_write/rgraynext[2] ), .CK(
        clk_30M), .RN(nReset), .Q(\fifo_write/rgray [2]) );
  DFFRHQ \fifo_write/wq1_rgray_reg[2]  ( .D(\fifo_write/rgray [2]), .CK(clk), 
        .RN(nReset), .Q(\fifo_write/wq1_rgray [2]) );
  DFFRHQ \fifo_write/wq2_rgray_reg[2]  ( .D(\fifo_write/wq1_rgray [2]), .CK(
        clk), .RN(nReset), .Q(\fifo_write/wq2_rgray [2]) );
  DFFRHQ \fifo_write/rbin_reg[4]  ( .D(\fifo_write/rbinnext[4] ), .CK(clk_30M), 
        .RN(nReset), .Q(\fifo_write/rbin[4] ) );
  DFFRHQ \fifo_write/rgray_reg[3]  ( .D(\fifo_write/rgraynext[3] ), .CK(
        clk_30M), .RN(nReset), .Q(\fifo_write/rgray [3]) );
  DFFRHQ \fifo_write/wq1_rgray_reg[3]  ( .D(\fifo_write/rgray [3]), .CK(clk), 
        .RN(nReset), .Q(\fifo_write/wq1_rgray [3]) );
  DFFRHQ \fifo_write/wq2_rgray_reg[3]  ( .D(\fifo_write/wq1_rgray [3]), .CK(
        clk), .RN(nReset), .Q(\fifo_write/wq2_rgray [3]) );
  DFFRHQ \fifo_write/rgray_reg[5]  ( .D(\fifo_write/rbinnext[5] ), .CK(clk_30M), .RN(nReset), .Q(\fifo_write/rgray [5]) );
  DFFRHQ \fifo_write/rgray_reg[4]  ( .D(\fifo_write/rgraynext[4] ), .CK(
        clk_30M), .RN(nReset), .Q(\fifo_write/rgray [4]) );
  DFFRHQ \fifo_write/wq1_rgray_reg[4]  ( .D(\fifo_write/rgray [4]), .CK(clk), 
        .RN(nReset), .Q(\fifo_write/wq1_rgray [4]) );
  DFFRHQ \fifo_write/wq2_rgray_reg[4]  ( .D(\fifo_write/wq1_rgray [4]), .CK(
        clk), .RN(nReset), .Q(\fifo_write/wq2_rgray [4]) );
  DFFHQ \fifo_write/mem_reg[16][7]  ( .D(n569), .CK(clk), .Q(
        \fifo_write/mem[16][7] ) );
  DFFHQ \fifo_write/mem_reg[16][6]  ( .D(n570), .CK(clk), .Q(
        \fifo_write/mem[16][6] ) );
  DFFHQ \fifo_write/mem_reg[16][5]  ( .D(n571), .CK(clk), .Q(
        \fifo_write/mem[16][5] ) );
  DFFHQ \fifo_write/mem_reg[16][4]  ( .D(n572), .CK(clk), .Q(
        \fifo_write/mem[16][4] ) );
  DFFHQ \fifo_write/mem_reg[16][3]  ( .D(n573), .CK(clk), .Q(
        \fifo_write/mem[16][3] ) );
  DFFHQ \fifo_write/mem_reg[16][2]  ( .D(n574), .CK(clk), .Q(
        \fifo_write/mem[16][2] ) );
  DFFHQ \fifo_write/mem_reg[16][1]  ( .D(n575), .CK(clk), .Q(
        \fifo_write/mem[16][1] ) );
  DFFHQ \fifo_write/mem_reg[16][0]  ( .D(n576), .CK(clk), .Q(
        \fifo_write/mem[16][0] ) );
  DFFHQ \fifo_write/mem_reg[17][7]  ( .D(n577), .CK(clk), .Q(
        \fifo_write/mem[17][7] ) );
  DFFHQ \fifo_write/mem_reg[17][6]  ( .D(n578), .CK(clk), .Q(
        \fifo_write/mem[17][6] ) );
  DFFHQ \fifo_write/mem_reg[17][5]  ( .D(n579), .CK(clk), .Q(
        \fifo_write/mem[17][5] ) );
  DFFHQ \fifo_write/mem_reg[17][4]  ( .D(n580), .CK(clk), .Q(
        \fifo_write/mem[17][4] ) );
  DFFHQ \fifo_write/mem_reg[17][3]  ( .D(n581), .CK(clk), .Q(
        \fifo_write/mem[17][3] ) );
  DFFHQ \fifo_write/mem_reg[17][2]  ( .D(n582), .CK(clk), .Q(
        \fifo_write/mem[17][2] ) );
  DFFHQ \fifo_write/mem_reg[17][1]  ( .D(n583), .CK(clk), .Q(
        \fifo_write/mem[17][1] ) );
  DFFHQ \fifo_write/mem_reg[17][0]  ( .D(n584), .CK(clk), .Q(
        \fifo_write/mem[17][0] ) );
  DFFHQ \fifo_write/mem_reg[18][7]  ( .D(n585), .CK(clk), .Q(
        \fifo_write/mem[18][7] ) );
  DFFHQ \fifo_write/mem_reg[18][6]  ( .D(n586), .CK(clk), .Q(
        \fifo_write/mem[18][6] ) );
  DFFHQ \fifo_write/mem_reg[18][5]  ( .D(n587), .CK(clk), .Q(
        \fifo_write/mem[18][5] ) );
  DFFHQ \fifo_write/mem_reg[18][4]  ( .D(n588), .CK(clk), .Q(
        \fifo_write/mem[18][4] ) );
  DFFHQ \fifo_write/mem_reg[18][3]  ( .D(n589), .CK(clk), .Q(
        \fifo_write/mem[18][3] ) );
  DFFHQ \fifo_write/mem_reg[18][2]  ( .D(n590), .CK(clk), .Q(
        \fifo_write/mem[18][2] ) );
  DFFHQ \fifo_write/mem_reg[18][1]  ( .D(n591), .CK(clk), .Q(
        \fifo_write/mem[18][1] ) );
  DFFHQ \fifo_write/mem_reg[18][0]  ( .D(n592), .CK(clk), .Q(
        \fifo_write/mem[18][0] ) );
  DFFHQ \fifo_write/mem_reg[19][7]  ( .D(n593), .CK(clk), .Q(
        \fifo_write/mem[19][7] ) );
  DFFHQ \fifo_write/mem_reg[19][6]  ( .D(n594), .CK(clk), .Q(
        \fifo_write/mem[19][6] ) );
  DFFHQ \fifo_write/mem_reg[19][5]  ( .D(n595), .CK(clk), .Q(
        \fifo_write/mem[19][5] ) );
  DFFHQ \fifo_write/mem_reg[19][4]  ( .D(n596), .CK(clk), .Q(
        \fifo_write/mem[19][4] ) );
  DFFHQ \fifo_write/mem_reg[19][3]  ( .D(n597), .CK(clk), .Q(
        \fifo_write/mem[19][3] ) );
  DFFHQ \fifo_write/mem_reg[19][2]  ( .D(n598), .CK(clk), .Q(
        \fifo_write/mem[19][2] ) );
  DFFHQ \fifo_write/mem_reg[19][1]  ( .D(n599), .CK(clk), .Q(
        \fifo_write/mem[19][1] ) );
  DFFHQ \fifo_write/mem_reg[19][0]  ( .D(n600), .CK(clk), .Q(
        \fifo_write/mem[19][0] ) );
  DFFHQ \fifo_write/mem_reg[20][7]  ( .D(n601), .CK(clk), .Q(
        \fifo_write/mem[20][7] ) );
  DFFHQ \fifo_write/mem_reg[20][6]  ( .D(n602), .CK(clk), .Q(
        \fifo_write/mem[20][6] ) );
  DFFHQ \fifo_write/mem_reg[20][5]  ( .D(n603), .CK(clk), .Q(
        \fifo_write/mem[20][5] ) );
  DFFHQ \fifo_write/mem_reg[20][4]  ( .D(n604), .CK(clk), .Q(
        \fifo_write/mem[20][4] ) );
  DFFHQ \fifo_write/mem_reg[20][3]  ( .D(n605), .CK(clk), .Q(
        \fifo_write/mem[20][3] ) );
  DFFHQ \fifo_write/mem_reg[20][2]  ( .D(n606), .CK(clk), .Q(
        \fifo_write/mem[20][2] ) );
  DFFHQ \fifo_write/mem_reg[20][1]  ( .D(n607), .CK(clk), .Q(
        \fifo_write/mem[20][1] ) );
  DFFHQ \fifo_write/mem_reg[20][0]  ( .D(n608), .CK(clk), .Q(
        \fifo_write/mem[20][0] ) );
  DFFHQ \fifo_write/mem_reg[21][7]  ( .D(n609), .CK(clk), .Q(
        \fifo_write/mem[21][7] ) );
  DFFHQ \fifo_write/mem_reg[21][6]  ( .D(n610), .CK(clk), .Q(
        \fifo_write/mem[21][6] ) );
  DFFHQ \fifo_write/mem_reg[21][5]  ( .D(n611), .CK(clk), .Q(
        \fifo_write/mem[21][5] ) );
  DFFHQ \fifo_write/mem_reg[21][4]  ( .D(n612), .CK(clk), .Q(
        \fifo_write/mem[21][4] ) );
  DFFHQ \fifo_write/mem_reg[21][3]  ( .D(n613), .CK(clk), .Q(
        \fifo_write/mem[21][3] ) );
  DFFHQ \fifo_write/mem_reg[21][2]  ( .D(n614), .CK(clk), .Q(
        \fifo_write/mem[21][2] ) );
  DFFHQ \fifo_write/mem_reg[21][1]  ( .D(n615), .CK(clk), .Q(
        \fifo_write/mem[21][1] ) );
  DFFHQ \fifo_write/mem_reg[21][0]  ( .D(n616), .CK(clk), .Q(
        \fifo_write/mem[21][0] ) );
  DFFHQ \fifo_write/mem_reg[22][7]  ( .D(n617), .CK(clk), .Q(
        \fifo_write/mem[22][7] ) );
  DFFHQ \fifo_write/mem_reg[22][6]  ( .D(n618), .CK(clk), .Q(
        \fifo_write/mem[22][6] ) );
  DFFHQ \fifo_write/mem_reg[22][5]  ( .D(n619), .CK(clk), .Q(
        \fifo_write/mem[22][5] ) );
  DFFHQ \fifo_write/mem_reg[22][4]  ( .D(n620), .CK(clk), .Q(
        \fifo_write/mem[22][4] ) );
  DFFHQ \fifo_write/mem_reg[22][3]  ( .D(n621), .CK(clk), .Q(
        \fifo_write/mem[22][3] ) );
  DFFHQ \fifo_write/mem_reg[22][2]  ( .D(n622), .CK(clk), .Q(
        \fifo_write/mem[22][2] ) );
  DFFHQ \fifo_write/mem_reg[22][1]  ( .D(n623), .CK(clk), .Q(
        \fifo_write/mem[22][1] ) );
  DFFHQ \fifo_write/mem_reg[22][0]  ( .D(n624), .CK(clk), .Q(
        \fifo_write/mem[22][0] ) );
  DFFHQ \fifo_write/mem_reg[23][7]  ( .D(n625), .CK(clk), .Q(
        \fifo_write/mem[23][7] ) );
  DFFHQ \fifo_write/mem_reg[23][6]  ( .D(n626), .CK(clk), .Q(
        \fifo_write/mem[23][6] ) );
  DFFHQ \fifo_write/mem_reg[23][5]  ( .D(n627), .CK(clk), .Q(
        \fifo_write/mem[23][5] ) );
  DFFHQ \fifo_write/mem_reg[23][4]  ( .D(n628), .CK(clk), .Q(
        \fifo_write/mem[23][4] ) );
  DFFHQ \fifo_write/mem_reg[23][3]  ( .D(n629), .CK(clk), .Q(
        \fifo_write/mem[23][3] ) );
  DFFHQ \fifo_write/mem_reg[23][2]  ( .D(n630), .CK(clk), .Q(
        \fifo_write/mem[23][2] ) );
  DFFHQ \fifo_write/mem_reg[23][1]  ( .D(n631), .CK(clk), .Q(
        \fifo_write/mem[23][1] ) );
  DFFHQ \fifo_write/mem_reg[23][0]  ( .D(n632), .CK(clk), .Q(
        \fifo_write/mem[23][0] ) );
  DFFHQ \fifo_write/mem_reg[0][7]  ( .D(n441), .CK(clk), .Q(
        \fifo_write/mem[0][7] ) );
  DFFHQ \fifo_write/mem_reg[0][6]  ( .D(n442), .CK(clk), .Q(
        \fifo_write/mem[0][6] ) );
  DFFHQ \fifo_write/mem_reg[0][5]  ( .D(n443), .CK(clk), .Q(
        \fifo_write/mem[0][5] ) );
  DFFHQ \fifo_write/mem_reg[0][4]  ( .D(n444), .CK(clk), .Q(
        \fifo_write/mem[0][4] ) );
  DFFHQ \fifo_write/mem_reg[0][3]  ( .D(n445), .CK(clk), .Q(
        \fifo_write/mem[0][3] ) );
  DFFHQ \fifo_write/mem_reg[0][2]  ( .D(n446), .CK(clk), .Q(
        \fifo_write/mem[0][2] ) );
  DFFHQ \fifo_write/mem_reg[0][1]  ( .D(n447), .CK(clk), .Q(
        \fifo_write/mem[0][1] ) );
  DFFHQ \fifo_write/mem_reg[0][0]  ( .D(n448), .CK(clk), .Q(
        \fifo_write/mem[0][0] ) );
  DFFHQ \fifo_write/mem_reg[1][7]  ( .D(n449), .CK(clk), .Q(
        \fifo_write/mem[1][7] ) );
  DFFHQ \fifo_write/mem_reg[1][6]  ( .D(n450), .CK(clk), .Q(
        \fifo_write/mem[1][6] ) );
  DFFHQ \fifo_write/mem_reg[1][5]  ( .D(n451), .CK(clk), .Q(
        \fifo_write/mem[1][5] ) );
  DFFHQ \fifo_write/mem_reg[1][4]  ( .D(n452), .CK(clk), .Q(
        \fifo_write/mem[1][4] ) );
  DFFHQ \fifo_write/mem_reg[1][3]  ( .D(n453), .CK(clk), .Q(
        \fifo_write/mem[1][3] ) );
  DFFHQ \fifo_write/mem_reg[1][2]  ( .D(n454), .CK(clk), .Q(
        \fifo_write/mem[1][2] ) );
  DFFHQ \fifo_write/mem_reg[1][1]  ( .D(n455), .CK(clk), .Q(
        \fifo_write/mem[1][1] ) );
  DFFHQ \fifo_write/mem_reg[1][0]  ( .D(n456), .CK(clk), .Q(
        \fifo_write/mem[1][0] ) );
  DFFHQ \fifo_write/mem_reg[2][7]  ( .D(n457), .CK(clk), .Q(
        \fifo_write/mem[2][7] ) );
  DFFHQ \fifo_write/mem_reg[2][6]  ( .D(n458), .CK(clk), .Q(
        \fifo_write/mem[2][6] ) );
  DFFHQ \fifo_write/mem_reg[2][5]  ( .D(n459), .CK(clk), .Q(
        \fifo_write/mem[2][5] ) );
  DFFHQ \fifo_write/mem_reg[2][4]  ( .D(n460), .CK(clk), .Q(
        \fifo_write/mem[2][4] ) );
  DFFHQ \fifo_write/mem_reg[2][3]  ( .D(n461), .CK(clk), .Q(
        \fifo_write/mem[2][3] ) );
  DFFHQ \fifo_write/mem_reg[2][2]  ( .D(n462), .CK(clk), .Q(
        \fifo_write/mem[2][2] ) );
  DFFHQ \fifo_write/mem_reg[2][1]  ( .D(n463), .CK(clk), .Q(
        \fifo_write/mem[2][1] ) );
  DFFHQ \fifo_write/mem_reg[2][0]  ( .D(n464), .CK(clk), .Q(
        \fifo_write/mem[2][0] ) );
  DFFHQ \fifo_write/mem_reg[3][7]  ( .D(n465), .CK(clk), .Q(
        \fifo_write/mem[3][7] ) );
  DFFHQ \fifo_write/mem_reg[3][6]  ( .D(n466), .CK(clk), .Q(
        \fifo_write/mem[3][6] ) );
  DFFHQ \fifo_write/mem_reg[3][5]  ( .D(n467), .CK(clk), .Q(
        \fifo_write/mem[3][5] ) );
  DFFHQ \fifo_write/mem_reg[3][4]  ( .D(n468), .CK(clk), .Q(
        \fifo_write/mem[3][4] ) );
  DFFHQ \fifo_write/mem_reg[3][3]  ( .D(n469), .CK(clk), .Q(
        \fifo_write/mem[3][3] ) );
  DFFHQ \fifo_write/mem_reg[3][2]  ( .D(n470), .CK(clk), .Q(
        \fifo_write/mem[3][2] ) );
  DFFHQ \fifo_write/mem_reg[3][1]  ( .D(n471), .CK(clk), .Q(
        \fifo_write/mem[3][1] ) );
  DFFHQ \fifo_write/mem_reg[3][0]  ( .D(n472), .CK(clk), .Q(
        \fifo_write/mem[3][0] ) );
  DFFHQ \fifo_write/mem_reg[4][7]  ( .D(n473), .CK(clk), .Q(
        \fifo_write/mem[4][7] ) );
  DFFHQ \fifo_write/mem_reg[4][6]  ( .D(n474), .CK(clk), .Q(
        \fifo_write/mem[4][6] ) );
  DFFHQ \fifo_write/mem_reg[4][5]  ( .D(n475), .CK(clk), .Q(
        \fifo_write/mem[4][5] ) );
  DFFHQ \fifo_write/mem_reg[4][4]  ( .D(n476), .CK(clk), .Q(
        \fifo_write/mem[4][4] ) );
  DFFHQ \fifo_write/mem_reg[4][3]  ( .D(n477), .CK(clk), .Q(
        \fifo_write/mem[4][3] ) );
  DFFHQ \fifo_write/mem_reg[4][2]  ( .D(n478), .CK(clk), .Q(
        \fifo_write/mem[4][2] ) );
  DFFHQ \fifo_write/mem_reg[4][1]  ( .D(n479), .CK(clk), .Q(
        \fifo_write/mem[4][1] ) );
  DFFHQ \fifo_write/mem_reg[4][0]  ( .D(n480), .CK(clk), .Q(
        \fifo_write/mem[4][0] ) );
  DFFHQ \fifo_write/mem_reg[5][7]  ( .D(n481), .CK(clk), .Q(
        \fifo_write/mem[5][7] ) );
  DFFHQ \fifo_write/mem_reg[5][6]  ( .D(n482), .CK(clk), .Q(
        \fifo_write/mem[5][6] ) );
  DFFHQ \fifo_write/mem_reg[5][5]  ( .D(n483), .CK(clk), .Q(
        \fifo_write/mem[5][5] ) );
  DFFHQ \fifo_write/mem_reg[5][4]  ( .D(n484), .CK(clk), .Q(
        \fifo_write/mem[5][4] ) );
  DFFHQ \fifo_write/mem_reg[5][3]  ( .D(n485), .CK(clk), .Q(
        \fifo_write/mem[5][3] ) );
  DFFHQ \fifo_write/mem_reg[5][2]  ( .D(n486), .CK(clk), .Q(
        \fifo_write/mem[5][2] ) );
  DFFHQ \fifo_write/mem_reg[5][1]  ( .D(n487), .CK(clk), .Q(
        \fifo_write/mem[5][1] ) );
  DFFHQ \fifo_write/mem_reg[5][0]  ( .D(n488), .CK(clk), .Q(
        \fifo_write/mem[5][0] ) );
  DFFHQ \fifo_write/mem_reg[6][7]  ( .D(n489), .CK(clk), .Q(
        \fifo_write/mem[6][7] ) );
  DFFHQ \fifo_write/mem_reg[6][6]  ( .D(n490), .CK(clk), .Q(
        \fifo_write/mem[6][6] ) );
  DFFHQ \fifo_write/mem_reg[6][5]  ( .D(n491), .CK(clk), .Q(
        \fifo_write/mem[6][5] ) );
  DFFHQ \fifo_write/mem_reg[6][4]  ( .D(n492), .CK(clk), .Q(
        \fifo_write/mem[6][4] ) );
  DFFHQ \fifo_write/mem_reg[6][3]  ( .D(n493), .CK(clk), .Q(
        \fifo_write/mem[6][3] ) );
  DFFHQ \fifo_write/mem_reg[6][2]  ( .D(n494), .CK(clk), .Q(
        \fifo_write/mem[6][2] ) );
  DFFHQ \fifo_write/mem_reg[6][1]  ( .D(n495), .CK(clk), .Q(
        \fifo_write/mem[6][1] ) );
  DFFHQ \fifo_write/mem_reg[6][0]  ( .D(n496), .CK(clk), .Q(
        \fifo_write/mem[6][0] ) );
  DFFHQ \fifo_write/mem_reg[7][7]  ( .D(n497), .CK(clk), .Q(
        \fifo_write/mem[7][7] ) );
  DFFHQ \fifo_write/mem_reg[7][6]  ( .D(n498), .CK(clk), .Q(
        \fifo_write/mem[7][6] ) );
  DFFHQ \fifo_write/mem_reg[7][5]  ( .D(n499), .CK(clk), .Q(
        \fifo_write/mem[7][5] ) );
  DFFHQ \fifo_write/mem_reg[7][4]  ( .D(n500), .CK(clk), .Q(
        \fifo_write/mem[7][4] ) );
  DFFHQ \fifo_write/mem_reg[7][3]  ( .D(n501), .CK(clk), .Q(
        \fifo_write/mem[7][3] ) );
  DFFHQ \fifo_write/mem_reg[7][2]  ( .D(n502), .CK(clk), .Q(
        \fifo_write/mem[7][2] ) );
  DFFHQ \fifo_write/mem_reg[7][1]  ( .D(n503), .CK(clk), .Q(
        \fifo_write/mem[7][1] ) );
  DFFHQ \fifo_write/mem_reg[7][0]  ( .D(n504), .CK(clk), .Q(
        \fifo_write/mem[7][0] ) );
  DFFHQ \fifo_write/mem_reg[8][7]  ( .D(n505), .CK(clk), .Q(
        \fifo_write/mem[8][7] ) );
  DFFHQ \fifo_write/mem_reg[8][6]  ( .D(n506), .CK(clk), .Q(
        \fifo_write/mem[8][6] ) );
  DFFHQ \fifo_write/mem_reg[8][5]  ( .D(n507), .CK(clk), .Q(
        \fifo_write/mem[8][5] ) );
  DFFHQ \fifo_write/mem_reg[8][4]  ( .D(n508), .CK(clk), .Q(
        \fifo_write/mem[8][4] ) );
  DFFHQ \fifo_write/mem_reg[8][3]  ( .D(n509), .CK(clk), .Q(
        \fifo_write/mem[8][3] ) );
  DFFHQ \fifo_write/mem_reg[8][2]  ( .D(n510), .CK(clk), .Q(
        \fifo_write/mem[8][2] ) );
  DFFHQ \fifo_write/mem_reg[8][1]  ( .D(n511), .CK(clk), .Q(
        \fifo_write/mem[8][1] ) );
  DFFHQ \fifo_write/mem_reg[8][0]  ( .D(n512), .CK(clk), .Q(
        \fifo_write/mem[8][0] ) );
  DFFHQ \fifo_write/mem_reg[9][7]  ( .D(n513), .CK(clk), .Q(
        \fifo_write/mem[9][7] ) );
  DFFHQ \fifo_write/mem_reg[9][6]  ( .D(n514), .CK(clk), .Q(
        \fifo_write/mem[9][6] ) );
  DFFHQ \fifo_write/mem_reg[9][5]  ( .D(n515), .CK(clk), .Q(
        \fifo_write/mem[9][5] ) );
  DFFHQ \fifo_write/mem_reg[9][4]  ( .D(n516), .CK(clk), .Q(
        \fifo_write/mem[9][4] ) );
  DFFHQ \fifo_write/mem_reg[9][3]  ( .D(n517), .CK(clk), .Q(
        \fifo_write/mem[9][3] ) );
  DFFHQ \fifo_write/mem_reg[9][2]  ( .D(n518), .CK(clk), .Q(
        \fifo_write/mem[9][2] ) );
  DFFHQ \fifo_write/mem_reg[9][1]  ( .D(n519), .CK(clk), .Q(
        \fifo_write/mem[9][1] ) );
  DFFHQ \fifo_write/mem_reg[9][0]  ( .D(n520), .CK(clk), .Q(
        \fifo_write/mem[9][0] ) );
  DFFHQ \fifo_write/mem_reg[10][7]  ( .D(n521), .CK(clk), .Q(
        \fifo_write/mem[10][7] ) );
  DFFHQ \fifo_write/mem_reg[10][6]  ( .D(n522), .CK(clk), .Q(
        \fifo_write/mem[10][6] ) );
  DFFHQ \fifo_write/mem_reg[10][5]  ( .D(n523), .CK(clk), .Q(
        \fifo_write/mem[10][5] ) );
  DFFHQ \fifo_write/mem_reg[10][4]  ( .D(n524), .CK(clk), .Q(
        \fifo_write/mem[10][4] ) );
  DFFHQ \fifo_write/mem_reg[10][3]  ( .D(n525), .CK(clk), .Q(
        \fifo_write/mem[10][3] ) );
  DFFHQ \fifo_write/mem_reg[10][2]  ( .D(n526), .CK(clk), .Q(
        \fifo_write/mem[10][2] ) );
  DFFHQ \fifo_write/mem_reg[10][1]  ( .D(n527), .CK(clk), .Q(
        \fifo_write/mem[10][1] ) );
  DFFHQ \fifo_write/mem_reg[10][0]  ( .D(n528), .CK(clk), .Q(
        \fifo_write/mem[10][0] ) );
  DFFHQ \fifo_write/mem_reg[11][7]  ( .D(n529), .CK(clk), .Q(
        \fifo_write/mem[11][7] ) );
  DFFHQ \fifo_write/mem_reg[11][6]  ( .D(n530), .CK(clk), .Q(
        \fifo_write/mem[11][6] ) );
  DFFHQ \fifo_write/mem_reg[11][5]  ( .D(n531), .CK(clk), .Q(
        \fifo_write/mem[11][5] ) );
  DFFHQ \fifo_write/mem_reg[11][4]  ( .D(n532), .CK(clk), .Q(
        \fifo_write/mem[11][4] ) );
  DFFHQ \fifo_write/mem_reg[11][3]  ( .D(n533), .CK(clk), .Q(
        \fifo_write/mem[11][3] ) );
  DFFHQ \fifo_write/mem_reg[11][2]  ( .D(n534), .CK(clk), .Q(
        \fifo_write/mem[11][2] ) );
  DFFHQ \fifo_write/mem_reg[11][1]  ( .D(n535), .CK(clk), .Q(
        \fifo_write/mem[11][1] ) );
  DFFHQ \fifo_write/mem_reg[11][0]  ( .D(n536), .CK(clk), .Q(
        \fifo_write/mem[11][0] ) );
  DFFHQ \fifo_write/mem_reg[12][7]  ( .D(n537), .CK(clk), .Q(
        \fifo_write/mem[12][7] ) );
  DFFHQ \fifo_write/mem_reg[12][6]  ( .D(n538), .CK(clk), .Q(
        \fifo_write/mem[12][6] ) );
  DFFHQ \fifo_write/mem_reg[12][5]  ( .D(n539), .CK(clk), .Q(
        \fifo_write/mem[12][5] ) );
  DFFHQ \fifo_write/mem_reg[12][4]  ( .D(n540), .CK(clk), .Q(
        \fifo_write/mem[12][4] ) );
  DFFHQ \fifo_write/mem_reg[12][3]  ( .D(n541), .CK(clk), .Q(
        \fifo_write/mem[12][3] ) );
  DFFHQ \fifo_write/mem_reg[12][2]  ( .D(n542), .CK(clk), .Q(
        \fifo_write/mem[12][2] ) );
  DFFHQ \fifo_write/mem_reg[12][1]  ( .D(n543), .CK(clk), .Q(
        \fifo_write/mem[12][1] ) );
  DFFHQ \fifo_write/mem_reg[12][0]  ( .D(n544), .CK(clk), .Q(
        \fifo_write/mem[12][0] ) );
  DFFHQ \fifo_write/mem_reg[13][7]  ( .D(n545), .CK(clk), .Q(
        \fifo_write/mem[13][7] ) );
  DFFHQ \fifo_write/mem_reg[13][6]  ( .D(n546), .CK(clk), .Q(
        \fifo_write/mem[13][6] ) );
  DFFHQ \fifo_write/mem_reg[13][5]  ( .D(n547), .CK(clk), .Q(
        \fifo_write/mem[13][5] ) );
  DFFHQ \fifo_write/mem_reg[13][4]  ( .D(n548), .CK(clk), .Q(
        \fifo_write/mem[13][4] ) );
  DFFHQ \fifo_write/mem_reg[13][3]  ( .D(n549), .CK(clk), .Q(
        \fifo_write/mem[13][3] ) );
  DFFHQ \fifo_write/mem_reg[13][2]  ( .D(n550), .CK(clk), .Q(
        \fifo_write/mem[13][2] ) );
  DFFHQ \fifo_write/mem_reg[13][1]  ( .D(n551), .CK(clk), .Q(
        \fifo_write/mem[13][1] ) );
  DFFHQ \fifo_write/mem_reg[13][0]  ( .D(n552), .CK(clk), .Q(
        \fifo_write/mem[13][0] ) );
  DFFHQ \fifo_write/mem_reg[14][7]  ( .D(n553), .CK(clk), .Q(
        \fifo_write/mem[14][7] ) );
  DFFHQ \fifo_write/mem_reg[14][6]  ( .D(n554), .CK(clk), .Q(
        \fifo_write/mem[14][6] ) );
  DFFHQ \fifo_write/mem_reg[14][5]  ( .D(n555), .CK(clk), .Q(
        \fifo_write/mem[14][5] ) );
  DFFHQ \fifo_write/mem_reg[14][4]  ( .D(n556), .CK(clk), .Q(
        \fifo_write/mem[14][4] ) );
  DFFHQ \fifo_write/mem_reg[14][3]  ( .D(n557), .CK(clk), .Q(
        \fifo_write/mem[14][3] ) );
  DFFHQ \fifo_write/mem_reg[14][2]  ( .D(n558), .CK(clk), .Q(
        \fifo_write/mem[14][2] ) );
  DFFHQ \fifo_write/mem_reg[14][1]  ( .D(n559), .CK(clk), .Q(
        \fifo_write/mem[14][1] ) );
  DFFHQ \fifo_write/mem_reg[14][0]  ( .D(n560), .CK(clk), .Q(
        \fifo_write/mem[14][0] ) );
  DFFHQ \fifo_write/mem_reg[15][7]  ( .D(n561), .CK(clk), .Q(
        \fifo_write/mem[15][7] ) );
  DFFHQ \fifo_write/mem_reg[15][6]  ( .D(n562), .CK(clk), .Q(
        \fifo_write/mem[15][6] ) );
  DFFHQ \fifo_write/mem_reg[15][5]  ( .D(n563), .CK(clk), .Q(
        \fifo_write/mem[15][5] ) );
  DFFHQ \fifo_write/mem_reg[15][4]  ( .D(n564), .CK(clk), .Q(
        \fifo_write/mem[15][4] ) );
  DFFHQ \fifo_write/mem_reg[15][3]  ( .D(n565), .CK(clk), .Q(
        \fifo_write/mem[15][3] ) );
  DFFHQ \fifo_write/mem_reg[15][2]  ( .D(n566), .CK(clk), .Q(
        \fifo_write/mem[15][2] ) );
  DFFHQ \fifo_write/mem_reg[15][1]  ( .D(n567), .CK(clk), .Q(
        \fifo_write/mem[15][1] ) );
  DFFHQ \fifo_write/mem_reg[15][0]  ( .D(n568), .CK(clk), .Q(
        \fifo_write/mem[15][0] ) );
  DFFHQ \fifo_write/mem_reg[24][7]  ( .D(n633), .CK(clk), .Q(
        \fifo_write/mem[24][7] ) );
  DFFHQ \fifo_write/mem_reg[24][6]  ( .D(n634), .CK(clk), .Q(
        \fifo_write/mem[24][6] ) );
  DFFHQ \fifo_write/mem_reg[24][5]  ( .D(n635), .CK(clk), .Q(
        \fifo_write/mem[24][5] ) );
  DFFHQ \fifo_write/mem_reg[24][4]  ( .D(n636), .CK(clk), .Q(
        \fifo_write/mem[24][4] ) );
  DFFHQ \fifo_write/mem_reg[24][3]  ( .D(n637), .CK(clk), .Q(
        \fifo_write/mem[24][3] ) );
  DFFHQ \fifo_write/mem_reg[24][2]  ( .D(n638), .CK(clk), .Q(
        \fifo_write/mem[24][2] ) );
  DFFHQ \fifo_write/mem_reg[24][1]  ( .D(n639), .CK(clk), .Q(
        \fifo_write/mem[24][1] ) );
  DFFHQ \fifo_write/mem_reg[24][0]  ( .D(n640), .CK(clk), .Q(
        \fifo_write/mem[24][0] ) );
  DFFHQ \fifo_write/mem_reg[25][7]  ( .D(n641), .CK(clk), .Q(
        \fifo_write/mem[25][7] ) );
  DFFHQ \fifo_write/mem_reg[25][6]  ( .D(n642), .CK(clk), .Q(
        \fifo_write/mem[25][6] ) );
  DFFHQ \fifo_write/mem_reg[25][5]  ( .D(n643), .CK(clk), .Q(
        \fifo_write/mem[25][5] ) );
  DFFHQ \fifo_write/mem_reg[25][4]  ( .D(n644), .CK(clk), .Q(
        \fifo_write/mem[25][4] ) );
  DFFHQ \fifo_write/mem_reg[25][3]  ( .D(n645), .CK(clk), .Q(
        \fifo_write/mem[25][3] ) );
  DFFHQ \fifo_write/mem_reg[25][2]  ( .D(n646), .CK(clk), .Q(
        \fifo_write/mem[25][2] ) );
  DFFHQ \fifo_write/mem_reg[25][1]  ( .D(n647), .CK(clk), .Q(
        \fifo_write/mem[25][1] ) );
  DFFHQ \fifo_write/mem_reg[25][0]  ( .D(n648), .CK(clk), .Q(
        \fifo_write/mem[25][0] ) );
  DFFHQ \fifo_write/mem_reg[26][7]  ( .D(n649), .CK(clk), .Q(
        \fifo_write/mem[26][7] ) );
  DFFHQ \fifo_write/mem_reg[26][6]  ( .D(n650), .CK(clk), .Q(
        \fifo_write/mem[26][6] ) );
  DFFHQ \fifo_write/mem_reg[26][5]  ( .D(n651), .CK(clk), .Q(
        \fifo_write/mem[26][5] ) );
  DFFHQ \fifo_write/mem_reg[26][4]  ( .D(n652), .CK(clk), .Q(
        \fifo_write/mem[26][4] ) );
  DFFHQ \fifo_write/mem_reg[26][3]  ( .D(n653), .CK(clk), .Q(
        \fifo_write/mem[26][3] ) );
  DFFHQ \fifo_write/mem_reg[26][2]  ( .D(n654), .CK(clk), .Q(
        \fifo_write/mem[26][2] ) );
  DFFHQ \fifo_write/mem_reg[26][1]  ( .D(n655), .CK(clk), .Q(
        \fifo_write/mem[26][1] ) );
  DFFHQ \fifo_write/mem_reg[26][0]  ( .D(n656), .CK(clk), .Q(
        \fifo_write/mem[26][0] ) );
  DFFHQ \fifo_write/mem_reg[27][7]  ( .D(n657), .CK(clk), .Q(
        \fifo_write/mem[27][7] ) );
  DFFHQ \fifo_write/mem_reg[27][6]  ( .D(n658), .CK(clk), .Q(
        \fifo_write/mem[27][6] ) );
  DFFHQ \fifo_write/mem_reg[27][5]  ( .D(n659), .CK(clk), .Q(
        \fifo_write/mem[27][5] ) );
  DFFHQ \fifo_write/mem_reg[27][4]  ( .D(n660), .CK(clk), .Q(
        \fifo_write/mem[27][4] ) );
  DFFHQ \fifo_write/mem_reg[27][3]  ( .D(n661), .CK(clk), .Q(
        \fifo_write/mem[27][3] ) );
  DFFHQ \fifo_write/mem_reg[27][2]  ( .D(n662), .CK(clk), .Q(
        \fifo_write/mem[27][2] ) );
  DFFHQ \fifo_write/mem_reg[27][1]  ( .D(n663), .CK(clk), .Q(
        \fifo_write/mem[27][1] ) );
  DFFHQ \fifo_write/mem_reg[27][0]  ( .D(n664), .CK(clk), .Q(
        \fifo_write/mem[27][0] ) );
  DFFHQ \fifo_write/mem_reg[28][7]  ( .D(n665), .CK(clk), .Q(
        \fifo_write/mem[28][7] ) );
  DFFHQ \fifo_write/mem_reg[28][6]  ( .D(n666), .CK(clk), .Q(
        \fifo_write/mem[28][6] ) );
  DFFHQ \fifo_write/mem_reg[28][5]  ( .D(n667), .CK(clk), .Q(
        \fifo_write/mem[28][5] ) );
  DFFHQ \fifo_write/mem_reg[28][4]  ( .D(n668), .CK(clk), .Q(
        \fifo_write/mem[28][4] ) );
  DFFHQ \fifo_write/mem_reg[28][3]  ( .D(n669), .CK(clk), .Q(
        \fifo_write/mem[28][3] ) );
  DFFHQ \fifo_write/mem_reg[28][2]  ( .D(n670), .CK(clk), .Q(
        \fifo_write/mem[28][2] ) );
  DFFHQ \fifo_write/mem_reg[28][1]  ( .D(n671), .CK(clk), .Q(
        \fifo_write/mem[28][1] ) );
  DFFHQ \fifo_write/mem_reg[28][0]  ( .D(n672), .CK(clk), .Q(
        \fifo_write/mem[28][0] ) );
  DFFHQ \fifo_write/mem_reg[29][7]  ( .D(n673), .CK(clk), .Q(
        \fifo_write/mem[29][7] ) );
  DFFHQ \fifo_write/mem_reg[29][6]  ( .D(n674), .CK(clk), .Q(
        \fifo_write/mem[29][6] ) );
  DFFHQ \fifo_write/mem_reg[29][5]  ( .D(n675), .CK(clk), .Q(
        \fifo_write/mem[29][5] ) );
  DFFHQ \fifo_write/mem_reg[29][4]  ( .D(n676), .CK(clk), .Q(
        \fifo_write/mem[29][4] ) );
  DFFHQ \fifo_write/mem_reg[29][3]  ( .D(n677), .CK(clk), .Q(
        \fifo_write/mem[29][3] ) );
  DFFHQ \fifo_write/mem_reg[29][2]  ( .D(n678), .CK(clk), .Q(
        \fifo_write/mem[29][2] ) );
  DFFHQ \fifo_write/mem_reg[29][1]  ( .D(n679), .CK(clk), .Q(
        \fifo_write/mem[29][1] ) );
  DFFHQ \fifo_write/mem_reg[29][0]  ( .D(n680), .CK(clk), .Q(
        \fifo_write/mem[29][0] ) );
  DFFHQ \fifo_write/mem_reg[30][7]  ( .D(n681), .CK(clk), .Q(
        \fifo_write/mem[30][7] ) );
  DFFHQ \fifo_write/mem_reg[30][6]  ( .D(n682), .CK(clk), .Q(
        \fifo_write/mem[30][6] ) );
  DFFHQ \fifo_write/mem_reg[30][5]  ( .D(n683), .CK(clk), .Q(
        \fifo_write/mem[30][5] ) );
  DFFHQ \fifo_write/mem_reg[30][4]  ( .D(n684), .CK(clk), .Q(
        \fifo_write/mem[30][4] ) );
  DFFHQ \fifo_write/mem_reg[30][3]  ( .D(n685), .CK(clk), .Q(
        \fifo_write/mem[30][3] ) );
  DFFHQ \fifo_write/mem_reg[30][2]  ( .D(n686), .CK(clk), .Q(
        \fifo_write/mem[30][2] ) );
  DFFHQ \fifo_write/mem_reg[30][1]  ( .D(n687), .CK(clk), .Q(
        \fifo_write/mem[30][1] ) );
  DFFHQ \fifo_write/mem_reg[30][0]  ( .D(n688), .CK(clk), .Q(
        \fifo_write/mem[30][0] ) );
  DFFHQ \fifo_write/mem_reg[31][7]  ( .D(n689), .CK(clk), .Q(
        \fifo_write/mem[31][7] ) );
  DFFHQ \fifo_write/mem_reg[31][6]  ( .D(n690), .CK(clk), .Q(
        \fifo_write/mem[31][6] ) );
  DFFHQ \fifo_write/mem_reg[31][5]  ( .D(n691), .CK(clk), .Q(
        \fifo_write/mem[31][5] ) );
  DFFHQ \fifo_write/mem_reg[31][4]  ( .D(n692), .CK(clk), .Q(
        \fifo_write/mem[31][4] ) );
  DFFHQ \fifo_write/mem_reg[31][3]  ( .D(n693), .CK(clk), .Q(
        \fifo_write/mem[31][3] ) );
  DFFHQ \fifo_write/mem_reg[31][2]  ( .D(n694), .CK(clk), .Q(
        \fifo_write/mem[31][2] ) );
  DFFHQ \fifo_write/mem_reg[31][1]  ( .D(n695), .CK(clk), .Q(
        \fifo_write/mem[31][1] ) );
  DFFHQ \fifo_write/mem_reg[31][0]  ( .D(n696), .CK(clk), .Q(
        \fifo_write/mem[31][0] ) );
  DFFRHQ \fifo_read/wq1_rgray_reg[5]  ( .D(\fifo_read/rgray [5]), .CK(clk_30M), 
        .RN(nReset), .Q(\fifo_read/wq1_rgray [5]) );
  DFFRHQ \fifo_read/wq2_rgray_reg[5]  ( .D(\fifo_read/wq1_rgray [5]), .CK(
        clk_30M), .RN(nReset), .Q(\fifo_read/wq2_rgray [5]) );
  DFFRHQ \fifo_read/o_wfull_reg  ( .D(\fifo_read/wfull_next ), .CK(clk_30M), 
        .RN(nReset), .Q(o_wfull) );
  DFFRHQ \fifo_read/wbin_reg[0]  ( .D(\fifo_read/wbinnext[0] ), .CK(clk_30M), 
        .RN(nReset), .Q(\fifo_read/waddr[0] ) );
  DFFRHQ \fifo_read/wbin_reg[1]  ( .D(\fifo_read/wbinnext[1] ), .CK(clk_30M), 
        .RN(nReset), .Q(\fifo_read/waddr[1] ) );
  DFFRHQ \fifo_read/wgray_reg[0]  ( .D(\fifo_read/wgraynext[0] ), .CK(clk_30M), 
        .RN(nReset), .Q(\fifo_read/wgray [0]) );
  DFFRHQ \fifo_read/rq1_wgray_reg[0]  ( .D(\fifo_read/wgray [0]), .CK(clk), 
        .RN(nReset), .Q(\fifo_read/rq1_wgray [0]) );
  DFFRHQ \fifo_read/rq2_wgray_reg[0]  ( .D(\fifo_read/rq1_wgray [0]), .CK(clk), 
        .RN(nReset), .Q(\fifo_read/rq2_wgray [0]) );
  DFFRHQ \fifo_read/wbin_reg[2]  ( .D(\fifo_read/wbinnext[2] ), .CK(clk_30M), 
        .RN(nReset), .Q(\fifo_read/waddr[2] ) );
  DFFRHQ \fifo_read/wgray_reg[1]  ( .D(\fifo_read/wgraynext[1] ), .CK(clk_30M), 
        .RN(nReset), .Q(\fifo_read/wgray [1]) );
  DFFRHQ \fifo_read/rq1_wgray_reg[1]  ( .D(\fifo_read/wgray [1]), .CK(clk), 
        .RN(nReset), .Q(\fifo_read/rq1_wgray [1]) );
  DFFRHQ \fifo_read/rq2_wgray_reg[1]  ( .D(\fifo_read/rq1_wgray [1]), .CK(clk), 
        .RN(nReset), .Q(\fifo_read/rq2_wgray [1]) );
  DFFRHQ \fifo_read/wbin_reg[3]  ( .D(\fifo_read/wbinnext[3] ), .CK(clk_30M), 
        .RN(nReset), .Q(\fifo_read/waddr[3] ) );
  DFFRHQ \fifo_read/wgray_reg[2]  ( .D(\fifo_read/wgraynext[2] ), .CK(clk_30M), 
        .RN(nReset), .Q(\fifo_read/wgray [2]) );
  DFFRHQ \fifo_read/rq1_wgray_reg[2]  ( .D(\fifo_read/wgray [2]), .CK(clk), 
        .RN(nReset), .Q(\fifo_read/rq1_wgray [2]) );
  DFFRHQ \fifo_read/rq2_wgray_reg[2]  ( .D(\fifo_read/rq1_wgray [2]), .CK(clk), 
        .RN(nReset), .Q(\fifo_read/rq2_wgray [2]) );
  DFFRHQ \fifo_read/wbin_reg[4]  ( .D(\fifo_read/wbinnext[4] ), .CK(clk_30M), 
        .RN(nReset), .Q(\fifo_read/waddr[4] ) );
  DFFRHQ \fifo_read/wgray_reg[3]  ( .D(\fifo_read/wgraynext[3] ), .CK(clk_30M), 
        .RN(nReset), .Q(\fifo_read/wgray [3]) );
  DFFRHQ \fifo_read/rq1_wgray_reg[3]  ( .D(\fifo_read/wgray [3]), .CK(clk), 
        .RN(nReset), .Q(\fifo_read/rq1_wgray [3]) );
  DFFRHQ \fifo_read/rq2_wgray_reg[3]  ( .D(\fifo_read/rq1_wgray [3]), .CK(clk), 
        .RN(nReset), .Q(\fifo_read/rq2_wgray [3]) );
  DFFRHQ \fifo_read/wgray_reg[5]  ( .D(\fifo_read/wbinnext[5] ), .CK(clk_30M), 
        .RN(nReset), .Q(\fifo_read/wgray [5]) );
  DFFRHQ \fifo_read/rq1_wgray_reg[5]  ( .D(\fifo_read/wgray [5]), .CK(clk), 
        .RN(nReset), .Q(\fifo_read/rq1_wgray [5]) );
  DFFRHQ \fifo_read/rq2_wgray_reg[5]  ( .D(\fifo_read/rq1_wgray [5]), .CK(clk), 
        .RN(nReset), .Q(\fifo_read/rq2_wgray [5]) );
  DFFRHQ \fifo_read/wgray_reg[4]  ( .D(\fifo_read/wgraynext[4] ), .CK(clk_30M), 
        .RN(nReset), .Q(\fifo_read/wgray [4]) );
  DFFRHQ \fifo_read/rq1_wgray_reg[4]  ( .D(\fifo_read/wgray [4]), .CK(clk), 
        .RN(nReset), .Q(\fifo_read/rq1_wgray [4]) );
  DFFRHQ \fifo_read/rq2_wgray_reg[4]  ( .D(\fifo_read/rq1_wgray [4]), .CK(clk), 
        .RN(nReset), .Q(\fifo_read/rq2_wgray [4]) );
  DFFSHQ \fifo_read/o_rempty_reg  ( .D(\fifo_read/rempty_next ), .CK(clk), 
        .SN(nReset), .Q(o_rempty) );
  DFFRHQ \fifo_read/rbin_reg[0]  ( .D(\fifo_read/rbinnext[0] ), .CK(clk), .RN(
        nReset), .Q(\fifo_read/rbin[0] ) );
  DFFRHQ \fifo_read/rbin_reg[1]  ( .D(\fifo_read/rbinnext[1] ), .CK(clk), .RN(
        nReset), .Q(\fifo_read/rbin[1] ) );
  DFFRHQ \fifo_read/rgray_reg[0]  ( .D(\fifo_read/rgraynext[0] ), .CK(clk), 
        .RN(nReset), .Q(\fifo_read/rgray [0]) );
  DFFRHQ \fifo_read/wq1_rgray_reg[0]  ( .D(\fifo_read/rgray [0]), .CK(clk_30M), 
        .RN(nReset), .Q(\fifo_read/wq1_rgray [0]) );
  DFFRHQ \fifo_read/wq2_rgray_reg[0]  ( .D(\fifo_read/wq1_rgray [0]), .CK(
        clk_30M), .RN(nReset), .Q(\fifo_read/wq2_rgray [0]) );
  DFFRHQ \fifo_read/rbin_reg[2]  ( .D(\fifo_read/rbinnext[2] ), .CK(clk), .RN(
        nReset), .Q(\fifo_read/rbin[2] ) );
  DFFRHQ \fifo_read/rgray_reg[1]  ( .D(\fifo_read/rgraynext[1] ), .CK(clk), 
        .RN(nReset), .Q(\fifo_read/rgray [1]) );
  DFFRHQ \fifo_read/wq1_rgray_reg[1]  ( .D(\fifo_read/rgray [1]), .CK(clk_30M), 
        .RN(nReset), .Q(\fifo_read/wq1_rgray [1]) );
  DFFRHQ \fifo_read/wq2_rgray_reg[1]  ( .D(\fifo_read/wq1_rgray [1]), .CK(
        clk_30M), .RN(nReset), .Q(\fifo_read/wq2_rgray [1]) );
  DFFRHQ \fifo_read/rbin_reg[3]  ( .D(\fifo_read/rbinnext[3] ), .CK(clk), .RN(
        nReset), .Q(\fifo_read/rbin[3] ) );
  DFFRHQ \fifo_read/rgray_reg[2]  ( .D(\fifo_read/rgraynext[2] ), .CK(clk), 
        .RN(nReset), .Q(\fifo_read/rgray [2]) );
  DFFRHQ \fifo_read/wq1_rgray_reg[2]  ( .D(\fifo_read/rgray [2]), .CK(clk_30M), 
        .RN(nReset), .Q(\fifo_read/wq1_rgray [2]) );
  DFFRHQ \fifo_read/wq2_rgray_reg[2]  ( .D(\fifo_read/wq1_rgray [2]), .CK(
        clk_30M), .RN(nReset), .Q(\fifo_read/wq2_rgray [2]) );
  DFFRHQ \fifo_read/rbin_reg[4]  ( .D(\fifo_read/rbinnext[4] ), .CK(clk), .RN(
        nReset), .Q(\fifo_read/rbin[4] ) );
  DFFRHQ \fifo_read/rgray_reg[3]  ( .D(\fifo_read/rgraynext[3] ), .CK(clk), 
        .RN(nReset), .Q(\fifo_read/rgray [3]) );
  DFFRHQ \fifo_read/wq1_rgray_reg[3]  ( .D(\fifo_read/rgray [3]), .CK(clk_30M), 
        .RN(nReset), .Q(\fifo_read/wq1_rgray [3]) );
  DFFRHQ \fifo_read/wq2_rgray_reg[3]  ( .D(\fifo_read/wq1_rgray [3]), .CK(
        clk_30M), .RN(nReset), .Q(\fifo_read/wq2_rgray [3]) );
  DFFRHQ \fifo_read/rgray_reg[5]  ( .D(\fifo_read/rbinnext[5] ), .CK(clk), 
        .RN(nReset), .Q(\fifo_read/rgray [5]) );
  DFFRHQ \fifo_read/rgray_reg[4]  ( .D(\fifo_read/rgraynext[4] ), .CK(clk), 
        .RN(nReset), .Q(\fifo_read/rgray [4]) );
  DFFRHQ \fifo_read/wq1_rgray_reg[4]  ( .D(\fifo_read/rgray [4]), .CK(clk_30M), 
        .RN(nReset), .Q(\fifo_read/wq1_rgray [4]) );
  DFFRHQ \fifo_read/wq2_rgray_reg[4]  ( .D(\fifo_read/wq1_rgray [4]), .CK(
        clk_30M), .RN(nReset), .Q(\fifo_read/wq2_rgray [4]) );
  DFFHQ \fifo_read/mem_reg[16][7]  ( .D(n313), .CK(clk_30M), .Q(
        \fifo_read/mem[16][7] ) );
  DFFHQ \fifo_read/mem_reg[16][6]  ( .D(n314), .CK(clk_30M), .Q(
        \fifo_read/mem[16][6] ) );
  DFFHQ \fifo_read/mem_reg[16][5]  ( .D(n315), .CK(clk_30M), .Q(
        \fifo_read/mem[16][5] ) );
  DFFHQ \fifo_read/mem_reg[16][4]  ( .D(n316), .CK(clk_30M), .Q(
        \fifo_read/mem[16][4] ) );
  DFFHQ \fifo_read/mem_reg[16][3]  ( .D(n317), .CK(clk_30M), .Q(
        \fifo_read/mem[16][3] ) );
  DFFHQ \fifo_read/mem_reg[16][2]  ( .D(n318), .CK(clk_30M), .Q(
        \fifo_read/mem[16][2] ) );
  DFFHQ \fifo_read/mem_reg[16][1]  ( .D(n319), .CK(clk_30M), .Q(
        \fifo_read/mem[16][1] ) );
  DFFHQ \fifo_read/mem_reg[16][0]  ( .D(n320), .CK(clk_30M), .Q(
        \fifo_read/mem[16][0] ) );
  DFFHQ \fifo_read/mem_reg[17][7]  ( .D(n321), .CK(clk_30M), .Q(
        \fifo_read/mem[17][7] ) );
  DFFHQ \fifo_read/mem_reg[17][6]  ( .D(n322), .CK(clk_30M), .Q(
        \fifo_read/mem[17][6] ) );
  DFFHQ \fifo_read/mem_reg[17][5]  ( .D(n323), .CK(clk_30M), .Q(
        \fifo_read/mem[17][5] ) );
  DFFHQ \fifo_read/mem_reg[17][4]  ( .D(n324), .CK(clk_30M), .Q(
        \fifo_read/mem[17][4] ) );
  DFFHQ \fifo_read/mem_reg[17][3]  ( .D(n325), .CK(clk_30M), .Q(
        \fifo_read/mem[17][3] ) );
  DFFHQ \fifo_read/mem_reg[17][2]  ( .D(n326), .CK(clk_30M), .Q(
        \fifo_read/mem[17][2] ) );
  DFFHQ \fifo_read/mem_reg[17][1]  ( .D(n327), .CK(clk_30M), .Q(
        \fifo_read/mem[17][1] ) );
  DFFHQ \fifo_read/mem_reg[17][0]  ( .D(n328), .CK(clk_30M), .Q(
        \fifo_read/mem[17][0] ) );
  DFFHQ \fifo_read/mem_reg[18][7]  ( .D(n329), .CK(clk_30M), .Q(
        \fifo_read/mem[18][7] ) );
  DFFHQ \fifo_read/mem_reg[18][6]  ( .D(n330), .CK(clk_30M), .Q(
        \fifo_read/mem[18][6] ) );
  DFFHQ \fifo_read/mem_reg[18][5]  ( .D(n331), .CK(clk_30M), .Q(
        \fifo_read/mem[18][5] ) );
  DFFHQ \fifo_read/mem_reg[18][4]  ( .D(n332), .CK(clk_30M), .Q(
        \fifo_read/mem[18][4] ) );
  DFFHQ \fifo_read/mem_reg[18][3]  ( .D(n333), .CK(clk_30M), .Q(
        \fifo_read/mem[18][3] ) );
  DFFHQ \fifo_read/mem_reg[18][2]  ( .D(n334), .CK(clk_30M), .Q(
        \fifo_read/mem[18][2] ) );
  DFFHQ \fifo_read/mem_reg[18][1]  ( .D(n335), .CK(clk_30M), .Q(
        \fifo_read/mem[18][1] ) );
  DFFHQ \fifo_read/mem_reg[18][0]  ( .D(n336), .CK(clk_30M), .Q(
        \fifo_read/mem[18][0] ) );
  DFFHQ \fifo_read/mem_reg[19][7]  ( .D(n337), .CK(clk_30M), .Q(
        \fifo_read/mem[19][7] ) );
  DFFHQ \fifo_read/mem_reg[19][6]  ( .D(n338), .CK(clk_30M), .Q(
        \fifo_read/mem[19][6] ) );
  DFFHQ \fifo_read/mem_reg[19][5]  ( .D(n339), .CK(clk_30M), .Q(
        \fifo_read/mem[19][5] ) );
  DFFHQ \fifo_read/mem_reg[19][4]  ( .D(n340), .CK(clk_30M), .Q(
        \fifo_read/mem[19][4] ) );
  DFFHQ \fifo_read/mem_reg[19][3]  ( .D(n341), .CK(clk_30M), .Q(
        \fifo_read/mem[19][3] ) );
  DFFHQ \fifo_read/mem_reg[19][2]  ( .D(n342), .CK(clk_30M), .Q(
        \fifo_read/mem[19][2] ) );
  DFFHQ \fifo_read/mem_reg[19][1]  ( .D(n343), .CK(clk_30M), .Q(
        \fifo_read/mem[19][1] ) );
  DFFHQ \fifo_read/mem_reg[19][0]  ( .D(n344), .CK(clk_30M), .Q(
        \fifo_read/mem[19][0] ) );
  DFFHQ \fifo_read/mem_reg[20][7]  ( .D(n345), .CK(clk_30M), .Q(
        \fifo_read/mem[20][7] ) );
  DFFHQ \fifo_read/mem_reg[20][6]  ( .D(n346), .CK(clk_30M), .Q(
        \fifo_read/mem[20][6] ) );
  DFFHQ \fifo_read/mem_reg[20][5]  ( .D(n347), .CK(clk_30M), .Q(
        \fifo_read/mem[20][5] ) );
  DFFHQ \fifo_read/mem_reg[20][4]  ( .D(n348), .CK(clk_30M), .Q(
        \fifo_read/mem[20][4] ) );
  DFFHQ \fifo_read/mem_reg[20][3]  ( .D(n349), .CK(clk_30M), .Q(
        \fifo_read/mem[20][3] ) );
  DFFHQ \fifo_read/mem_reg[20][2]  ( .D(n350), .CK(clk_30M), .Q(
        \fifo_read/mem[20][2] ) );
  DFFHQ \fifo_read/mem_reg[20][1]  ( .D(n351), .CK(clk_30M), .Q(
        \fifo_read/mem[20][1] ) );
  DFFHQ \fifo_read/mem_reg[20][0]  ( .D(n352), .CK(clk_30M), .Q(
        \fifo_read/mem[20][0] ) );
  DFFHQ \fifo_read/mem_reg[21][7]  ( .D(n353), .CK(clk_30M), .Q(
        \fifo_read/mem[21][7] ) );
  DFFHQ \fifo_read/mem_reg[21][6]  ( .D(n354), .CK(clk_30M), .Q(
        \fifo_read/mem[21][6] ) );
  DFFHQ \fifo_read/mem_reg[21][5]  ( .D(n355), .CK(clk_30M), .Q(
        \fifo_read/mem[21][5] ) );
  DFFHQ \fifo_read/mem_reg[21][4]  ( .D(n356), .CK(clk_30M), .Q(
        \fifo_read/mem[21][4] ) );
  DFFHQ \fifo_read/mem_reg[21][3]  ( .D(n357), .CK(clk_30M), .Q(
        \fifo_read/mem[21][3] ) );
  DFFHQ \fifo_read/mem_reg[21][2]  ( .D(n358), .CK(clk_30M), .Q(
        \fifo_read/mem[21][2] ) );
  DFFHQ \fifo_read/mem_reg[21][1]  ( .D(n359), .CK(clk_30M), .Q(
        \fifo_read/mem[21][1] ) );
  DFFHQ \fifo_read/mem_reg[21][0]  ( .D(n360), .CK(clk_30M), .Q(
        \fifo_read/mem[21][0] ) );
  DFFHQ \fifo_read/mem_reg[22][7]  ( .D(n361), .CK(clk_30M), .Q(
        \fifo_read/mem[22][7] ) );
  DFFHQ \fifo_read/mem_reg[22][6]  ( .D(n362), .CK(clk_30M), .Q(
        \fifo_read/mem[22][6] ) );
  DFFHQ \fifo_read/mem_reg[22][5]  ( .D(n363), .CK(clk_30M), .Q(
        \fifo_read/mem[22][5] ) );
  DFFHQ \fifo_read/mem_reg[22][4]  ( .D(n364), .CK(clk_30M), .Q(
        \fifo_read/mem[22][4] ) );
  DFFHQ \fifo_read/mem_reg[22][3]  ( .D(n365), .CK(clk_30M), .Q(
        \fifo_read/mem[22][3] ) );
  DFFHQ \fifo_read/mem_reg[22][2]  ( .D(n366), .CK(clk_30M), .Q(
        \fifo_read/mem[22][2] ) );
  DFFHQ \fifo_read/mem_reg[22][1]  ( .D(n367), .CK(clk_30M), .Q(
        \fifo_read/mem[22][1] ) );
  DFFHQ \fifo_read/mem_reg[22][0]  ( .D(n368), .CK(clk_30M), .Q(
        \fifo_read/mem[22][0] ) );
  DFFHQ \fifo_read/mem_reg[23][7]  ( .D(n369), .CK(clk_30M), .Q(
        \fifo_read/mem[23][7] ) );
  DFFHQ \fifo_read/mem_reg[23][6]  ( .D(n370), .CK(clk_30M), .Q(
        \fifo_read/mem[23][6] ) );
  DFFHQ \fifo_read/mem_reg[23][5]  ( .D(n371), .CK(clk_30M), .Q(
        \fifo_read/mem[23][5] ) );
  DFFHQ \fifo_read/mem_reg[23][4]  ( .D(n372), .CK(clk_30M), .Q(
        \fifo_read/mem[23][4] ) );
  DFFHQ \fifo_read/mem_reg[23][3]  ( .D(n373), .CK(clk_30M), .Q(
        \fifo_read/mem[23][3] ) );
  DFFHQ \fifo_read/mem_reg[23][2]  ( .D(n374), .CK(clk_30M), .Q(
        \fifo_read/mem[23][2] ) );
  DFFHQ \fifo_read/mem_reg[23][1]  ( .D(n375), .CK(clk_30M), .Q(
        \fifo_read/mem[23][1] ) );
  DFFHQ \fifo_read/mem_reg[23][0]  ( .D(n376), .CK(clk_30M), .Q(
        \fifo_read/mem[23][0] ) );
  DFFHQ \fifo_read/mem_reg[0][7]  ( .D(n185), .CK(clk_30M), .Q(
        \fifo_read/mem[0][7] ) );
  DFFHQ \fifo_read/mem_reg[0][6]  ( .D(n186), .CK(clk_30M), .Q(
        \fifo_read/mem[0][6] ) );
  DFFHQ \fifo_read/mem_reg[0][5]  ( .D(n187), .CK(clk_30M), .Q(
        \fifo_read/mem[0][5] ) );
  DFFHQ \fifo_read/mem_reg[0][4]  ( .D(n188), .CK(clk_30M), .Q(
        \fifo_read/mem[0][4] ) );
  DFFHQ \fifo_read/mem_reg[0][3]  ( .D(n189), .CK(clk_30M), .Q(
        \fifo_read/mem[0][3] ) );
  DFFHQ \fifo_read/mem_reg[0][2]  ( .D(n190), .CK(clk_30M), .Q(
        \fifo_read/mem[0][2] ) );
  DFFHQ \fifo_read/mem_reg[0][1]  ( .D(n191), .CK(clk_30M), .Q(
        \fifo_read/mem[0][1] ) );
  DFFHQ \fifo_read/mem_reg[0][0]  ( .D(n192), .CK(clk_30M), .Q(
        \fifo_read/mem[0][0] ) );
  DFFHQ \fifo_read/mem_reg[1][7]  ( .D(n193), .CK(clk_30M), .Q(
        \fifo_read/mem[1][7] ) );
  DFFHQ \fifo_read/mem_reg[1][6]  ( .D(n194), .CK(clk_30M), .Q(
        \fifo_read/mem[1][6] ) );
  DFFHQ \fifo_read/mem_reg[1][5]  ( .D(n195), .CK(clk_30M), .Q(
        \fifo_read/mem[1][5] ) );
  DFFHQ \fifo_read/mem_reg[1][4]  ( .D(n196), .CK(clk_30M), .Q(
        \fifo_read/mem[1][4] ) );
  DFFHQ \fifo_read/mem_reg[1][3]  ( .D(n197), .CK(clk_30M), .Q(
        \fifo_read/mem[1][3] ) );
  DFFHQ \fifo_read/mem_reg[1][2]  ( .D(n198), .CK(clk_30M), .Q(
        \fifo_read/mem[1][2] ) );
  DFFHQ \fifo_read/mem_reg[1][1]  ( .D(n199), .CK(clk_30M), .Q(
        \fifo_read/mem[1][1] ) );
  DFFHQ \fifo_read/mem_reg[1][0]  ( .D(n200), .CK(clk_30M), .Q(
        \fifo_read/mem[1][0] ) );
  DFFHQ \fifo_read/mem_reg[2][7]  ( .D(n201), .CK(clk_30M), .Q(
        \fifo_read/mem[2][7] ) );
  DFFHQ \fifo_read/mem_reg[2][6]  ( .D(n202), .CK(clk_30M), .Q(
        \fifo_read/mem[2][6] ) );
  DFFHQ \fifo_read/mem_reg[2][5]  ( .D(n203), .CK(clk_30M), .Q(
        \fifo_read/mem[2][5] ) );
  DFFHQ \fifo_read/mem_reg[2][4]  ( .D(n204), .CK(clk_30M), .Q(
        \fifo_read/mem[2][4] ) );
  DFFHQ \fifo_read/mem_reg[2][3]  ( .D(n205), .CK(clk_30M), .Q(
        \fifo_read/mem[2][3] ) );
  DFFHQ \fifo_read/mem_reg[2][2]  ( .D(n206), .CK(clk_30M), .Q(
        \fifo_read/mem[2][2] ) );
  DFFHQ \fifo_read/mem_reg[2][1]  ( .D(n207), .CK(clk_30M), .Q(
        \fifo_read/mem[2][1] ) );
  DFFHQ \fifo_read/mem_reg[2][0]  ( .D(n208), .CK(clk_30M), .Q(
        \fifo_read/mem[2][0] ) );
  DFFHQ \fifo_read/mem_reg[3][7]  ( .D(n209), .CK(clk_30M), .Q(
        \fifo_read/mem[3][7] ) );
  DFFHQ \fifo_read/mem_reg[3][6]  ( .D(n210), .CK(clk_30M), .Q(
        \fifo_read/mem[3][6] ) );
  DFFHQ \fifo_read/mem_reg[3][5]  ( .D(n211), .CK(clk_30M), .Q(
        \fifo_read/mem[3][5] ) );
  DFFHQ \fifo_read/mem_reg[3][4]  ( .D(n212), .CK(clk_30M), .Q(
        \fifo_read/mem[3][4] ) );
  DFFHQ \fifo_read/mem_reg[3][3]  ( .D(n213), .CK(clk_30M), .Q(
        \fifo_read/mem[3][3] ) );
  DFFHQ \fifo_read/mem_reg[3][2]  ( .D(n214), .CK(clk_30M), .Q(
        \fifo_read/mem[3][2] ) );
  DFFHQ \fifo_read/mem_reg[3][1]  ( .D(n215), .CK(clk_30M), .Q(
        \fifo_read/mem[3][1] ) );
  DFFHQ \fifo_read/mem_reg[3][0]  ( .D(n216), .CK(clk_30M), .Q(
        \fifo_read/mem[3][0] ) );
  DFFHQ \fifo_read/mem_reg[4][7]  ( .D(n217), .CK(clk_30M), .Q(
        \fifo_read/mem[4][7] ) );
  DFFHQ \fifo_read/mem_reg[4][6]  ( .D(n218), .CK(clk_30M), .Q(
        \fifo_read/mem[4][6] ) );
  DFFHQ \fifo_read/mem_reg[4][5]  ( .D(n219), .CK(clk_30M), .Q(
        \fifo_read/mem[4][5] ) );
  DFFHQ \fifo_read/mem_reg[4][4]  ( .D(n220), .CK(clk_30M), .Q(
        \fifo_read/mem[4][4] ) );
  DFFHQ \fifo_read/mem_reg[4][3]  ( .D(n221), .CK(clk_30M), .Q(
        \fifo_read/mem[4][3] ) );
  DFFHQ \fifo_read/mem_reg[4][2]  ( .D(n222), .CK(clk_30M), .Q(
        \fifo_read/mem[4][2] ) );
  DFFHQ \fifo_read/mem_reg[4][1]  ( .D(n223), .CK(clk_30M), .Q(
        \fifo_read/mem[4][1] ) );
  DFFHQ \fifo_read/mem_reg[4][0]  ( .D(n224), .CK(clk_30M), .Q(
        \fifo_read/mem[4][0] ) );
  DFFHQ \fifo_read/mem_reg[5][7]  ( .D(n225), .CK(clk_30M), .Q(
        \fifo_read/mem[5][7] ) );
  DFFHQ \fifo_read/mem_reg[5][6]  ( .D(n226), .CK(clk_30M), .Q(
        \fifo_read/mem[5][6] ) );
  DFFHQ \fifo_read/mem_reg[5][5]  ( .D(n227), .CK(clk_30M), .Q(
        \fifo_read/mem[5][5] ) );
  DFFHQ \fifo_read/mem_reg[5][4]  ( .D(n228), .CK(clk_30M), .Q(
        \fifo_read/mem[5][4] ) );
  DFFHQ \fifo_read/mem_reg[5][3]  ( .D(n229), .CK(clk_30M), .Q(
        \fifo_read/mem[5][3] ) );
  DFFHQ \fifo_read/mem_reg[5][2]  ( .D(n230), .CK(clk_30M), .Q(
        \fifo_read/mem[5][2] ) );
  DFFHQ \fifo_read/mem_reg[5][1]  ( .D(n231), .CK(clk_30M), .Q(
        \fifo_read/mem[5][1] ) );
  DFFHQ \fifo_read/mem_reg[5][0]  ( .D(n232), .CK(clk_30M), .Q(
        \fifo_read/mem[5][0] ) );
  DFFHQ \fifo_read/mem_reg[6][7]  ( .D(n233), .CK(clk_30M), .Q(
        \fifo_read/mem[6][7] ) );
  DFFHQ \fifo_read/mem_reg[6][6]  ( .D(n234), .CK(clk_30M), .Q(
        \fifo_read/mem[6][6] ) );
  DFFHQ \fifo_read/mem_reg[6][5]  ( .D(n235), .CK(clk_30M), .Q(
        \fifo_read/mem[6][5] ) );
  DFFHQ \fifo_read/mem_reg[6][4]  ( .D(n236), .CK(clk_30M), .Q(
        \fifo_read/mem[6][4] ) );
  DFFHQ \fifo_read/mem_reg[6][3]  ( .D(n237), .CK(clk_30M), .Q(
        \fifo_read/mem[6][3] ) );
  DFFHQ \fifo_read/mem_reg[6][2]  ( .D(n238), .CK(clk_30M), .Q(
        \fifo_read/mem[6][2] ) );
  DFFHQ \fifo_read/mem_reg[6][1]  ( .D(n239), .CK(clk_30M), .Q(
        \fifo_read/mem[6][1] ) );
  DFFHQ \fifo_read/mem_reg[6][0]  ( .D(n240), .CK(clk_30M), .Q(
        \fifo_read/mem[6][0] ) );
  DFFHQ \fifo_read/mem_reg[7][7]  ( .D(n241), .CK(clk_30M), .Q(
        \fifo_read/mem[7][7] ) );
  DFFHQ \fifo_read/mem_reg[7][6]  ( .D(n242), .CK(clk_30M), .Q(
        \fifo_read/mem[7][6] ) );
  DFFHQ \fifo_read/mem_reg[7][5]  ( .D(n243), .CK(clk_30M), .Q(
        \fifo_read/mem[7][5] ) );
  DFFHQ \fifo_read/mem_reg[7][4]  ( .D(n244), .CK(clk_30M), .Q(
        \fifo_read/mem[7][4] ) );
  DFFHQ \fifo_read/mem_reg[7][3]  ( .D(n245), .CK(clk_30M), .Q(
        \fifo_read/mem[7][3] ) );
  DFFHQ \fifo_read/mem_reg[7][2]  ( .D(n246), .CK(clk_30M), .Q(
        \fifo_read/mem[7][2] ) );
  DFFHQ \fifo_read/mem_reg[7][1]  ( .D(n247), .CK(clk_30M), .Q(
        \fifo_read/mem[7][1] ) );
  DFFHQ \fifo_read/mem_reg[7][0]  ( .D(n248), .CK(clk_30M), .Q(
        \fifo_read/mem[7][0] ) );
  DFFHQ \fifo_read/mem_reg[8][7]  ( .D(n249), .CK(clk_30M), .Q(
        \fifo_read/mem[8][7] ) );
  DFFHQ \fifo_read/mem_reg[8][6]  ( .D(n250), .CK(clk_30M), .Q(
        \fifo_read/mem[8][6] ) );
  DFFHQ \fifo_read/mem_reg[8][5]  ( .D(n251), .CK(clk_30M), .Q(
        \fifo_read/mem[8][5] ) );
  DFFHQ \fifo_read/mem_reg[8][4]  ( .D(n252), .CK(clk_30M), .Q(
        \fifo_read/mem[8][4] ) );
  DFFHQ \fifo_read/mem_reg[8][3]  ( .D(n253), .CK(clk_30M), .Q(
        \fifo_read/mem[8][3] ) );
  DFFHQ \fifo_read/mem_reg[8][2]  ( .D(n254), .CK(clk_30M), .Q(
        \fifo_read/mem[8][2] ) );
  DFFHQ \fifo_read/mem_reg[8][1]  ( .D(n255), .CK(clk_30M), .Q(
        \fifo_read/mem[8][1] ) );
  DFFHQ \fifo_read/mem_reg[8][0]  ( .D(n256), .CK(clk_30M), .Q(
        \fifo_read/mem[8][0] ) );
  DFFHQ \fifo_read/mem_reg[9][7]  ( .D(n257), .CK(clk_30M), .Q(
        \fifo_read/mem[9][7] ) );
  DFFHQ \fifo_read/mem_reg[9][6]  ( .D(n258), .CK(clk_30M), .Q(
        \fifo_read/mem[9][6] ) );
  DFFHQ \fifo_read/mem_reg[9][5]  ( .D(n259), .CK(clk_30M), .Q(
        \fifo_read/mem[9][5] ) );
  DFFHQ \fifo_read/mem_reg[9][4]  ( .D(n260), .CK(clk_30M), .Q(
        \fifo_read/mem[9][4] ) );
  DFFHQ \fifo_read/mem_reg[9][3]  ( .D(n261), .CK(clk_30M), .Q(
        \fifo_read/mem[9][3] ) );
  DFFHQ \fifo_read/mem_reg[9][2]  ( .D(n262), .CK(clk_30M), .Q(
        \fifo_read/mem[9][2] ) );
  DFFHQ \fifo_read/mem_reg[9][1]  ( .D(n263), .CK(clk_30M), .Q(
        \fifo_read/mem[9][1] ) );
  DFFHQ \fifo_read/mem_reg[9][0]  ( .D(n264), .CK(clk_30M), .Q(
        \fifo_read/mem[9][0] ) );
  DFFHQ \fifo_read/mem_reg[10][7]  ( .D(n265), .CK(clk_30M), .Q(
        \fifo_read/mem[10][7] ) );
  DFFHQ \fifo_read/mem_reg[10][6]  ( .D(n266), .CK(clk_30M), .Q(
        \fifo_read/mem[10][6] ) );
  DFFHQ \fifo_read/mem_reg[10][5]  ( .D(n267), .CK(clk_30M), .Q(
        \fifo_read/mem[10][5] ) );
  DFFHQ \fifo_read/mem_reg[10][4]  ( .D(n268), .CK(clk_30M), .Q(
        \fifo_read/mem[10][4] ) );
  DFFHQ \fifo_read/mem_reg[10][3]  ( .D(n269), .CK(clk_30M), .Q(
        \fifo_read/mem[10][3] ) );
  DFFHQ \fifo_read/mem_reg[10][2]  ( .D(n270), .CK(clk_30M), .Q(
        \fifo_read/mem[10][2] ) );
  DFFHQ \fifo_read/mem_reg[10][1]  ( .D(n271), .CK(clk_30M), .Q(
        \fifo_read/mem[10][1] ) );
  DFFHQ \fifo_read/mem_reg[10][0]  ( .D(n272), .CK(clk_30M), .Q(
        \fifo_read/mem[10][0] ) );
  DFFHQ \fifo_read/mem_reg[11][7]  ( .D(n273), .CK(clk_30M), .Q(
        \fifo_read/mem[11][7] ) );
  DFFHQ \fifo_read/mem_reg[11][6]  ( .D(n274), .CK(clk_30M), .Q(
        \fifo_read/mem[11][6] ) );
  DFFHQ \fifo_read/mem_reg[11][5]  ( .D(n275), .CK(clk_30M), .Q(
        \fifo_read/mem[11][5] ) );
  DFFHQ \fifo_read/mem_reg[11][4]  ( .D(n276), .CK(clk_30M), .Q(
        \fifo_read/mem[11][4] ) );
  DFFHQ \fifo_read/mem_reg[11][3]  ( .D(n277), .CK(clk_30M), .Q(
        \fifo_read/mem[11][3] ) );
  DFFHQ \fifo_read/mem_reg[11][2]  ( .D(n278), .CK(clk_30M), .Q(
        \fifo_read/mem[11][2] ) );
  DFFHQ \fifo_read/mem_reg[11][1]  ( .D(n279), .CK(clk_30M), .Q(
        \fifo_read/mem[11][1] ) );
  DFFHQ \fifo_read/mem_reg[11][0]  ( .D(n280), .CK(clk_30M), .Q(
        \fifo_read/mem[11][0] ) );
  DFFHQ \fifo_read/mem_reg[12][7]  ( .D(n281), .CK(clk_30M), .Q(
        \fifo_read/mem[12][7] ) );
  DFFHQ \fifo_read/mem_reg[12][6]  ( .D(n282), .CK(clk_30M), .Q(
        \fifo_read/mem[12][6] ) );
  DFFHQ \fifo_read/mem_reg[12][5]  ( .D(n283), .CK(clk_30M), .Q(
        \fifo_read/mem[12][5] ) );
  DFFHQ \fifo_read/mem_reg[12][4]  ( .D(n284), .CK(clk_30M), .Q(
        \fifo_read/mem[12][4] ) );
  DFFHQ \fifo_read/mem_reg[12][3]  ( .D(n285), .CK(clk_30M), .Q(
        \fifo_read/mem[12][3] ) );
  DFFHQ \fifo_read/mem_reg[12][2]  ( .D(n286), .CK(clk_30M), .Q(
        \fifo_read/mem[12][2] ) );
  DFFHQ \fifo_read/mem_reg[12][1]  ( .D(n287), .CK(clk_30M), .Q(
        \fifo_read/mem[12][1] ) );
  DFFHQ \fifo_read/mem_reg[12][0]  ( .D(n288), .CK(clk_30M), .Q(
        \fifo_read/mem[12][0] ) );
  DFFHQ \fifo_read/mem_reg[13][7]  ( .D(n289), .CK(clk_30M), .Q(
        \fifo_read/mem[13][7] ) );
  DFFHQ \fifo_read/mem_reg[13][6]  ( .D(n290), .CK(clk_30M), .Q(
        \fifo_read/mem[13][6] ) );
  DFFHQ \fifo_read/mem_reg[13][5]  ( .D(n291), .CK(clk_30M), .Q(
        \fifo_read/mem[13][5] ) );
  DFFHQ \fifo_read/mem_reg[13][4]  ( .D(n292), .CK(clk_30M), .Q(
        \fifo_read/mem[13][4] ) );
  DFFHQ \fifo_read/mem_reg[13][3]  ( .D(n293), .CK(clk_30M), .Q(
        \fifo_read/mem[13][3] ) );
  DFFHQ \fifo_read/mem_reg[13][2]  ( .D(n294), .CK(clk_30M), .Q(
        \fifo_read/mem[13][2] ) );
  DFFHQ \fifo_read/mem_reg[13][1]  ( .D(n295), .CK(clk_30M), .Q(
        \fifo_read/mem[13][1] ) );
  DFFHQ \fifo_read/mem_reg[13][0]  ( .D(n296), .CK(clk_30M), .Q(
        \fifo_read/mem[13][0] ) );
  DFFHQ \fifo_read/mem_reg[14][7]  ( .D(n297), .CK(clk_30M), .Q(
        \fifo_read/mem[14][7] ) );
  DFFHQ \fifo_read/mem_reg[14][6]  ( .D(n298), .CK(clk_30M), .Q(
        \fifo_read/mem[14][6] ) );
  DFFHQ \fifo_read/mem_reg[14][5]  ( .D(n299), .CK(clk_30M), .Q(
        \fifo_read/mem[14][5] ) );
  DFFHQ \fifo_read/mem_reg[14][4]  ( .D(n300), .CK(clk_30M), .Q(
        \fifo_read/mem[14][4] ) );
  DFFHQ \fifo_read/mem_reg[14][3]  ( .D(n301), .CK(clk_30M), .Q(
        \fifo_read/mem[14][3] ) );
  DFFHQ \fifo_read/mem_reg[14][2]  ( .D(n302), .CK(clk_30M), .Q(
        \fifo_read/mem[14][2] ) );
  DFFHQ \fifo_read/mem_reg[14][1]  ( .D(n303), .CK(clk_30M), .Q(
        \fifo_read/mem[14][1] ) );
  DFFHQ \fifo_read/mem_reg[14][0]  ( .D(n304), .CK(clk_30M), .Q(
        \fifo_read/mem[14][0] ) );
  DFFHQ \fifo_read/mem_reg[15][7]  ( .D(n305), .CK(clk_30M), .Q(
        \fifo_read/mem[15][7] ) );
  DFFHQ \fifo_read/mem_reg[15][6]  ( .D(n306), .CK(clk_30M), .Q(
        \fifo_read/mem[15][6] ) );
  DFFHQ \fifo_read/mem_reg[15][5]  ( .D(n307), .CK(clk_30M), .Q(
        \fifo_read/mem[15][5] ) );
  DFFHQ \fifo_read/mem_reg[15][4]  ( .D(n308), .CK(clk_30M), .Q(
        \fifo_read/mem[15][4] ) );
  DFFHQ \fifo_read/mem_reg[15][3]  ( .D(n309), .CK(clk_30M), .Q(
        \fifo_read/mem[15][3] ) );
  DFFHQ \fifo_read/mem_reg[15][2]  ( .D(n310), .CK(clk_30M), .Q(
        \fifo_read/mem[15][2] ) );
  DFFHQ \fifo_read/mem_reg[15][1]  ( .D(n311), .CK(clk_30M), .Q(
        \fifo_read/mem[15][1] ) );
  DFFHQ \fifo_read/mem_reg[15][0]  ( .D(n312), .CK(clk_30M), .Q(
        \fifo_read/mem[15][0] ) );
  DFFHQ \fifo_read/mem_reg[24][7]  ( .D(n377), .CK(clk_30M), .Q(
        \fifo_read/mem[24][7] ) );
  DFFHQ \fifo_read/mem_reg[24][6]  ( .D(n378), .CK(clk_30M), .Q(
        \fifo_read/mem[24][6] ) );
  DFFHQ \fifo_read/mem_reg[24][5]  ( .D(n379), .CK(clk_30M), .Q(
        \fifo_read/mem[24][5] ) );
  DFFHQ \fifo_read/mem_reg[24][4]  ( .D(n380), .CK(clk_30M), .Q(
        \fifo_read/mem[24][4] ) );
  DFFHQ \fifo_read/mem_reg[24][3]  ( .D(n381), .CK(clk_30M), .Q(
        \fifo_read/mem[24][3] ) );
  DFFHQ \fifo_read/mem_reg[24][2]  ( .D(n382), .CK(clk_30M), .Q(
        \fifo_read/mem[24][2] ) );
  DFFHQ \fifo_read/mem_reg[24][1]  ( .D(n383), .CK(clk_30M), .Q(
        \fifo_read/mem[24][1] ) );
  DFFHQ \fifo_read/mem_reg[24][0]  ( .D(n384), .CK(clk_30M), .Q(
        \fifo_read/mem[24][0] ) );
  DFFHQ \fifo_read/mem_reg[25][7]  ( .D(n385), .CK(clk_30M), .Q(
        \fifo_read/mem[25][7] ) );
  DFFHQ \fifo_read/mem_reg[25][6]  ( .D(n386), .CK(clk_30M), .Q(
        \fifo_read/mem[25][6] ) );
  DFFHQ \fifo_read/mem_reg[25][5]  ( .D(n387), .CK(clk_30M), .Q(
        \fifo_read/mem[25][5] ) );
  DFFHQ \fifo_read/mem_reg[25][4]  ( .D(n388), .CK(clk_30M), .Q(
        \fifo_read/mem[25][4] ) );
  DFFHQ \fifo_read/mem_reg[25][3]  ( .D(n389), .CK(clk_30M), .Q(
        \fifo_read/mem[25][3] ) );
  DFFHQ \fifo_read/mem_reg[25][2]  ( .D(n390), .CK(clk_30M), .Q(
        \fifo_read/mem[25][2] ) );
  DFFHQ \fifo_read/mem_reg[25][1]  ( .D(n391), .CK(clk_30M), .Q(
        \fifo_read/mem[25][1] ) );
  DFFHQ \fifo_read/mem_reg[25][0]  ( .D(n392), .CK(clk_30M), .Q(
        \fifo_read/mem[25][0] ) );
  DFFHQ \fifo_read/mem_reg[26][7]  ( .D(n393), .CK(clk_30M), .Q(
        \fifo_read/mem[26][7] ) );
  DFFHQ \fifo_read/mem_reg[26][6]  ( .D(n394), .CK(clk_30M), .Q(
        \fifo_read/mem[26][6] ) );
  DFFHQ \fifo_read/mem_reg[26][5]  ( .D(n395), .CK(clk_30M), .Q(
        \fifo_read/mem[26][5] ) );
  DFFHQ \fifo_read/mem_reg[26][4]  ( .D(n396), .CK(clk_30M), .Q(
        \fifo_read/mem[26][4] ) );
  DFFHQ \fifo_read/mem_reg[26][3]  ( .D(n397), .CK(clk_30M), .Q(
        \fifo_read/mem[26][3] ) );
  DFFHQ \fifo_read/mem_reg[26][2]  ( .D(n398), .CK(clk_30M), .Q(
        \fifo_read/mem[26][2] ) );
  DFFHQ \fifo_read/mem_reg[26][1]  ( .D(n399), .CK(clk_30M), .Q(
        \fifo_read/mem[26][1] ) );
  DFFHQ \fifo_read/mem_reg[26][0]  ( .D(n400), .CK(clk_30M), .Q(
        \fifo_read/mem[26][0] ) );
  DFFHQ \fifo_read/mem_reg[27][7]  ( .D(n401), .CK(clk_30M), .Q(
        \fifo_read/mem[27][7] ) );
  DFFHQ \fifo_read/mem_reg[27][6]  ( .D(n402), .CK(clk_30M), .Q(
        \fifo_read/mem[27][6] ) );
  DFFHQ \fifo_read/mem_reg[27][5]  ( .D(n403), .CK(clk_30M), .Q(
        \fifo_read/mem[27][5] ) );
  DFFHQ \fifo_read/mem_reg[27][4]  ( .D(n404), .CK(clk_30M), .Q(
        \fifo_read/mem[27][4] ) );
  DFFHQ \fifo_read/mem_reg[27][3]  ( .D(n405), .CK(clk_30M), .Q(
        \fifo_read/mem[27][3] ) );
  DFFHQ \fifo_read/mem_reg[27][2]  ( .D(n406), .CK(clk_30M), .Q(
        \fifo_read/mem[27][2] ) );
  DFFHQ \fifo_read/mem_reg[27][1]  ( .D(n407), .CK(clk_30M), .Q(
        \fifo_read/mem[27][1] ) );
  DFFHQ \fifo_read/mem_reg[27][0]  ( .D(n408), .CK(clk_30M), .Q(
        \fifo_read/mem[27][0] ) );
  DFFHQ \fifo_read/mem_reg[28][7]  ( .D(n409), .CK(clk_30M), .Q(
        \fifo_read/mem[28][7] ) );
  DFFHQ \fifo_read/mem_reg[28][6]  ( .D(n410), .CK(clk_30M), .Q(
        \fifo_read/mem[28][6] ) );
  DFFHQ \fifo_read/mem_reg[28][5]  ( .D(n411), .CK(clk_30M), .Q(
        \fifo_read/mem[28][5] ) );
  DFFHQ \fifo_read/mem_reg[28][4]  ( .D(n412), .CK(clk_30M), .Q(
        \fifo_read/mem[28][4] ) );
  DFFHQ \fifo_read/mem_reg[28][3]  ( .D(n413), .CK(clk_30M), .Q(
        \fifo_read/mem[28][3] ) );
  DFFHQ \fifo_read/mem_reg[28][2]  ( .D(n414), .CK(clk_30M), .Q(
        \fifo_read/mem[28][2] ) );
  DFFHQ \fifo_read/mem_reg[28][1]  ( .D(n415), .CK(clk_30M), .Q(
        \fifo_read/mem[28][1] ) );
  DFFHQ \fifo_read/mem_reg[28][0]  ( .D(n416), .CK(clk_30M), .Q(
        \fifo_read/mem[28][0] ) );
  DFFHQ \fifo_read/mem_reg[29][7]  ( .D(n417), .CK(clk_30M), .Q(
        \fifo_read/mem[29][7] ) );
  DFFHQ \fifo_read/mem_reg[29][6]  ( .D(n418), .CK(clk_30M), .Q(
        \fifo_read/mem[29][6] ) );
  DFFHQ \fifo_read/mem_reg[29][5]  ( .D(n419), .CK(clk_30M), .Q(
        \fifo_read/mem[29][5] ) );
  DFFHQ \fifo_read/mem_reg[29][4]  ( .D(n420), .CK(clk_30M), .Q(
        \fifo_read/mem[29][4] ) );
  DFFHQ \fifo_read/mem_reg[29][3]  ( .D(n421), .CK(clk_30M), .Q(
        \fifo_read/mem[29][3] ) );
  DFFHQ \fifo_read/mem_reg[29][2]  ( .D(n422), .CK(clk_30M), .Q(
        \fifo_read/mem[29][2] ) );
  DFFHQ \fifo_read/mem_reg[29][1]  ( .D(n423), .CK(clk_30M), .Q(
        \fifo_read/mem[29][1] ) );
  DFFHQ \fifo_read/mem_reg[29][0]  ( .D(n424), .CK(clk_30M), .Q(
        \fifo_read/mem[29][0] ) );
  DFFHQ \fifo_read/mem_reg[30][7]  ( .D(n425), .CK(clk_30M), .Q(
        \fifo_read/mem[30][7] ) );
  DFFHQ \fifo_read/mem_reg[30][6]  ( .D(n426), .CK(clk_30M), .Q(
        \fifo_read/mem[30][6] ) );
  DFFHQ \fifo_read/mem_reg[30][5]  ( .D(n427), .CK(clk_30M), .Q(
        \fifo_read/mem[30][5] ) );
  DFFHQ \fifo_read/mem_reg[30][4]  ( .D(n428), .CK(clk_30M), .Q(
        \fifo_read/mem[30][4] ) );
  DFFHQ \fifo_read/mem_reg[30][3]  ( .D(n429), .CK(clk_30M), .Q(
        \fifo_read/mem[30][3] ) );
  DFFHQ \fifo_read/mem_reg[30][2]  ( .D(n430), .CK(clk_30M), .Q(
        \fifo_read/mem[30][2] ) );
  DFFHQ \fifo_read/mem_reg[30][1]  ( .D(n431), .CK(clk_30M), .Q(
        \fifo_read/mem[30][1] ) );
  DFFHQ \fifo_read/mem_reg[30][0]  ( .D(n432), .CK(clk_30M), .Q(
        \fifo_read/mem[30][0] ) );
  DFFHQ \fifo_read/mem_reg[31][7]  ( .D(n433), .CK(clk_30M), .Q(
        \fifo_read/mem[31][7] ) );
  DFFHQ \fifo_read/mem_reg[31][6]  ( .D(n434), .CK(clk_30M), .Q(
        \fifo_read/mem[31][6] ) );
  DFFHQ \fifo_read/mem_reg[31][5]  ( .D(n435), .CK(clk_30M), .Q(
        \fifo_read/mem[31][5] ) );
  DFFHQ \fifo_read/mem_reg[31][4]  ( .D(n436), .CK(clk_30M), .Q(
        \fifo_read/mem[31][4] ) );
  DFFHQ \fifo_read/mem_reg[31][3]  ( .D(n437), .CK(clk_30M), .Q(
        \fifo_read/mem[31][3] ) );
  DFFHQ \fifo_read/mem_reg[31][2]  ( .D(n438), .CK(clk_30M), .Q(
        \fifo_read/mem[31][2] ) );
  DFFHQ \fifo_read/mem_reg[31][1]  ( .D(n439), .CK(clk_30M), .Q(
        \fifo_read/mem[31][1] ) );
  DFFHQ \fifo_read/mem_reg[31][0]  ( .D(n440), .CK(clk_30M), .Q(
        \fifo_read/mem[31][0] ) );
  MX2 U728 ( .A(\fifo_write/mem[0][0] ), .B(\fifo_write/mem[1][0] ), .S0(n1361), .Y(n697) );
  MX2 U729 ( .A(\fifo_write/mem[2][0] ), .B(\fifo_write/mem[3][0] ), .S0(n1367), .Y(n698) );
  MX2 U730 ( .A(\fifo_write/mem[4][0] ), .B(\fifo_write/mem[5][0] ), .S0(n1363), .Y(n699) );
  MX2 U731 ( .A(\fifo_write/mem[6][0] ), .B(\fifo_write/mem[7][0] ), .S0(n1359), .Y(n700) );
  MX2 U732 ( .A(\fifo_write/mem[8][0] ), .B(\fifo_write/mem[9][0] ), .S0(n1361), .Y(n701) );
  MX2 U733 ( .A(\fifo_write/mem[10][0] ), .B(\fifo_write/mem[11][0] ), .S0(
        n1359), .Y(n702) );
  MX2 U734 ( .A(\fifo_write/mem[12][0] ), .B(\fifo_write/mem[13][0] ), .S0(
        n1366), .Y(n703) );
  MX2 U735 ( .A(\fifo_write/mem[14][0] ), .B(\fifo_write/mem[15][0] ), .S0(
        n1365), .Y(n704) );
  MX2 U736 ( .A(\fifo_write/mem[16][0] ), .B(\fifo_write/mem[17][0] ), .S0(
        n1364), .Y(n705) );
  MX2 U737 ( .A(\fifo_write/mem[18][0] ), .B(\fifo_write/mem[19][0] ), .S0(
        n1362), .Y(n706) );
  MX2 U738 ( .A(\fifo_write/mem[20][0] ), .B(\fifo_write/mem[21][0] ), .S0(
        n1359), .Y(n707) );
  MX2 U739 ( .A(\fifo_write/mem[22][0] ), .B(\fifo_write/mem[23][0] ), .S0(
        n1360), .Y(n708) );
  MX2 U740 ( .A(\fifo_write/mem[24][0] ), .B(\fifo_write/mem[25][0] ), .S0(
        n1361), .Y(n709) );
  MX2 U741 ( .A(\fifo_write/mem[26][0] ), .B(\fifo_write/mem[27][0] ), .S0(
        n1367), .Y(n710) );
  MX2 U742 ( .A(\fifo_write/mem[28][0] ), .B(\fifo_write/mem[29][0] ), .S0(
        n1367), .Y(n711) );
  MX2 U743 ( .A(\fifo_write/mem[30][0] ), .B(\fifo_write/mem[31][0] ), .S0(
        n1367), .Y(n712) );
  MX2 U744 ( .A(n697), .B(n698), .S0(n1184), .Y(n713) );
  MX2 U745 ( .A(n699), .B(n700), .S0(n1342), .Y(n714) );
  MX2 U746 ( .A(n701), .B(n702), .S0(n1342), .Y(n715) );
  MX2 U747 ( .A(n703), .B(n704), .S0(n1341), .Y(n716) );
  MX2 U748 ( .A(n705), .B(n706), .S0(n1183), .Y(n717) );
  MX2 U749 ( .A(n707), .B(n708), .S0(n1342), .Y(n718) );
  MX2 U750 ( .A(n709), .B(n710), .S0(n1342), .Y(n719) );
  MX2 U751 ( .A(n711), .B(n712), .S0(n1342), .Y(n720) );
  MX2 U752 ( .A(n713), .B(n714), .S0(n1347), .Y(n721) );
  MX2 U753 ( .A(n715), .B(n716), .S0(\fifo_write/rbin[2] ), .Y(n722) );
  MX2 U754 ( .A(n717), .B(n718), .S0(n1348), .Y(n723) );
  MX2 U755 ( .A(n719), .B(n720), .S0(n1347), .Y(n724) );
  MX2 U756 ( .A(n721), .B(n722), .S0(\fifo_write/rbin[3] ), .Y(n725) );
  MX2 U757 ( .A(n723), .B(n724), .S0(n1332), .Y(n726) );
  MX2 U758 ( .A(n725), .B(n726), .S0(n1188), .Y(wdata_to_fifo[0]) );
  MX2 U759 ( .A(\fifo_write/mem[0][1] ), .B(\fifo_write/mem[1][1] ), .S0(n1367), .Y(n727) );
  MX2 U760 ( .A(\fifo_write/mem[2][1] ), .B(\fifo_write/mem[3][1] ), .S0(
        \fifo_write/rbin[0] ), .Y(n728) );
  MX2 U761 ( .A(\fifo_write/mem[4][1] ), .B(\fifo_write/mem[5][1] ), .S0(n1367), .Y(n729) );
  MX2 U762 ( .A(\fifo_write/mem[6][1] ), .B(\fifo_write/mem[7][1] ), .S0(
        \fifo_write/rbin[0] ), .Y(n730) );
  MX2 U763 ( .A(\fifo_write/mem[8][1] ), .B(\fifo_write/mem[9][1] ), .S0(n1367), .Y(n731) );
  MX2 U764 ( .A(\fifo_write/mem[10][1] ), .B(\fifo_write/mem[11][1] ), .S0(
        \fifo_write/rbin[0] ), .Y(n732) );
  MX2 U765 ( .A(\fifo_write/mem[12][1] ), .B(\fifo_write/mem[13][1] ), .S0(
        n1367), .Y(n733) );
  MX2 U766 ( .A(\fifo_write/mem[14][1] ), .B(\fifo_write/mem[15][1] ), .S0(
        \fifo_write/rbin[0] ), .Y(n734) );
  MX2 U767 ( .A(\fifo_write/mem[16][1] ), .B(\fifo_write/mem[17][1] ), .S0(
        n1367), .Y(n735) );
  MX2 U768 ( .A(\fifo_write/mem[18][1] ), .B(\fifo_write/mem[19][1] ), .S0(
        \fifo_write/rbin[0] ), .Y(n736) );
  MX2 U769 ( .A(\fifo_write/mem[20][1] ), .B(\fifo_write/mem[21][1] ), .S0(
        \fifo_write/rbin[0] ), .Y(n737) );
  MX2 U770 ( .A(\fifo_write/mem[22][1] ), .B(\fifo_write/mem[23][1] ), .S0(
        n1359), .Y(n738) );
  MX2 U771 ( .A(\fifo_write/mem[24][1] ), .B(\fifo_write/mem[25][1] ), .S0(
        n1359), .Y(n739) );
  MX2 U772 ( .A(\fifo_write/mem[26][1] ), .B(\fifo_write/mem[27][1] ), .S0(
        n1359), .Y(n740) );
  MX2 U773 ( .A(\fifo_write/mem[28][1] ), .B(\fifo_write/mem[29][1] ), .S0(
        n1359), .Y(n741) );
  MX2 U774 ( .A(\fifo_write/mem[30][1] ), .B(\fifo_write/mem[31][1] ), .S0(
        n1359), .Y(n742) );
  MX2 U775 ( .A(n727), .B(n728), .S0(n1184), .Y(n743) );
  MX2 U776 ( .A(n729), .B(n730), .S0(n1341), .Y(n744) );
  MX2 U777 ( .A(n731), .B(n732), .S0(n1341), .Y(n745) );
  MX2 U778 ( .A(n733), .B(n734), .S0(n1341), .Y(n746) );
  MX2 U779 ( .A(n735), .B(n736), .S0(n1183), .Y(n747) );
  MX2 U780 ( .A(n737), .B(n738), .S0(\fifo_write/rbin[1] ), .Y(n748) );
  MX2 U781 ( .A(n739), .B(n740), .S0(n1184), .Y(n749) );
  MX2 U782 ( .A(n741), .B(n742), .S0(n1184), .Y(n750) );
  MX2 U783 ( .A(n743), .B(n744), .S0(\fifo_write/rbin[2] ), .Y(n751) );
  MX2 U784 ( .A(n745), .B(n746), .S0(n1348), .Y(n752) );
  MX2 U785 ( .A(n747), .B(n748), .S0(n1347), .Y(n753) );
  MX2 U786 ( .A(n749), .B(n750), .S0(\fifo_write/rbin[2] ), .Y(n754) );
  MX2 U787 ( .A(n751), .B(n752), .S0(\fifo_write/rbin[3] ), .Y(n755) );
  MX2 U788 ( .A(n753), .B(n754), .S0(n1332), .Y(n756) );
  MX2 U789 ( .A(n755), .B(n756), .S0(n1188), .Y(wdata_to_fifo[1]) );
  MX2 U790 ( .A(\fifo_write/mem[0][2] ), .B(\fifo_write/mem[1][2] ), .S0(n1359), .Y(n757) );
  MX2 U791 ( .A(\fifo_write/mem[2][2] ), .B(\fifo_write/mem[3][2] ), .S0(n1359), .Y(n758) );
  MX2 U792 ( .A(\fifo_write/mem[4][2] ), .B(\fifo_write/mem[5][2] ), .S0(n1359), .Y(n759) );
  MX2 U793 ( .A(\fifo_write/mem[6][2] ), .B(\fifo_write/mem[7][2] ), .S0(n1359), .Y(n760) );
  MX2 U794 ( .A(\fifo_write/mem[8][2] ), .B(\fifo_write/mem[9][2] ), .S0(n1360), .Y(n761) );
  MX2 U795 ( .A(\fifo_write/mem[10][2] ), .B(\fifo_write/mem[11][2] ), .S0(
        n1360), .Y(n762) );
  MX2 U796 ( .A(\fifo_write/mem[12][2] ), .B(\fifo_write/mem[13][2] ), .S0(
        n1360), .Y(n763) );
  MX2 U797 ( .A(\fifo_write/mem[14][2] ), .B(\fifo_write/mem[15][2] ), .S0(
        n1360), .Y(n764) );
  MX2 U798 ( .A(\fifo_write/mem[16][2] ), .B(\fifo_write/mem[17][2] ), .S0(
        n1360), .Y(n765) );
  MX2 U799 ( .A(\fifo_write/mem[18][2] ), .B(\fifo_write/mem[19][2] ), .S0(
        n1360), .Y(n766) );
  MX2 U800 ( .A(\fifo_write/mem[20][2] ), .B(\fifo_write/mem[21][2] ), .S0(
        n1360), .Y(n767) );
  MX2 U801 ( .A(\fifo_write/mem[22][2] ), .B(\fifo_write/mem[23][2] ), .S0(
        n1360), .Y(n768) );
  MX2 U802 ( .A(\fifo_write/mem[24][2] ), .B(\fifo_write/mem[25][2] ), .S0(
        n1360), .Y(n769) );
  MX2 U803 ( .A(\fifo_write/mem[26][2] ), .B(\fifo_write/mem[27][2] ), .S0(
        n1361), .Y(n770) );
  MX2 U804 ( .A(\fifo_write/mem[28][2] ), .B(\fifo_write/mem[29][2] ), .S0(
        n1361), .Y(n771) );
  MX2 U805 ( .A(\fifo_write/mem[30][2] ), .B(\fifo_write/mem[31][2] ), .S0(
        n1361), .Y(n772) );
  MX2 U806 ( .A(n757), .B(n758), .S0(n1184), .Y(n773) );
  MX2 U807 ( .A(n759), .B(n760), .S0(n1183), .Y(n774) );
  MX2 U808 ( .A(n761), .B(n762), .S0(n1183), .Y(n775) );
  MX2 U809 ( .A(n763), .B(n764), .S0(n1184), .Y(n776) );
  MX2 U810 ( .A(n765), .B(n766), .S0(n1183), .Y(n777) );
  MX2 U811 ( .A(n767), .B(n768), .S0(n1342), .Y(n778) );
  MX2 U812 ( .A(n769), .B(n770), .S0(n1342), .Y(n779) );
  MX2 U813 ( .A(n771), .B(n772), .S0(n1342), .Y(n780) );
  MX2 U814 ( .A(n773), .B(n774), .S0(n1348), .Y(n781) );
  MX2 U815 ( .A(n775), .B(n776), .S0(n1347), .Y(n782) );
  MX2 U816 ( .A(n777), .B(n778), .S0(\fifo_write/rbin[2] ), .Y(n783) );
  MX2 U817 ( .A(n779), .B(n780), .S0(n1348), .Y(n784) );
  MX2 U818 ( .A(n781), .B(n782), .S0(\fifo_write/rbin[3] ), .Y(n785) );
  MX2 U819 ( .A(n783), .B(n784), .S0(n1332), .Y(n786) );
  MX2 U820 ( .A(n785), .B(n786), .S0(n1188), .Y(wdata_to_fifo[2]) );
  MX2 U821 ( .A(\fifo_write/mem[0][3] ), .B(\fifo_write/mem[1][3] ), .S0(n1361), .Y(n787) );
  MX2 U822 ( .A(\fifo_write/mem[2][3] ), .B(\fifo_write/mem[3][3] ), .S0(n1361), .Y(n788) );
  MX2 U823 ( .A(\fifo_write/mem[4][3] ), .B(\fifo_write/mem[5][3] ), .S0(n1361), .Y(n789) );
  MX2 U824 ( .A(\fifo_write/mem[6][3] ), .B(\fifo_write/mem[7][3] ), .S0(n1361), .Y(n790) );
  MX2 U825 ( .A(\fifo_write/mem[8][3] ), .B(\fifo_write/mem[9][3] ), .S0(n1361), .Y(n791) );
  MX2 U826 ( .A(\fifo_write/mem[10][3] ), .B(\fifo_write/mem[11][3] ), .S0(
        n1361), .Y(n792) );
  MX2 U827 ( .A(\fifo_write/mem[12][3] ), .B(\fifo_write/mem[13][3] ), .S0(
        n1362), .Y(n793) );
  MX2 U828 ( .A(\fifo_write/mem[14][3] ), .B(\fifo_write/mem[15][3] ), .S0(
        n1362), .Y(n794) );
  MX2 U829 ( .A(\fifo_write/mem[16][3] ), .B(\fifo_write/mem[17][3] ), .S0(
        n1362), .Y(n795) );
  MX2 U830 ( .A(\fifo_write/mem[18][3] ), .B(\fifo_write/mem[19][3] ), .S0(
        n1362), .Y(n796) );
  MX2 U831 ( .A(\fifo_write/mem[20][3] ), .B(\fifo_write/mem[21][3] ), .S0(
        n1362), .Y(n797) );
  MX2 U832 ( .A(\fifo_write/mem[22][3] ), .B(\fifo_write/mem[23][3] ), .S0(
        n1362), .Y(n798) );
  MX2 U833 ( .A(\fifo_write/mem[24][3] ), .B(\fifo_write/mem[25][3] ), .S0(
        n1362), .Y(n799) );
  MX2 U834 ( .A(\fifo_write/mem[26][3] ), .B(\fifo_write/mem[27][3] ), .S0(
        n1362), .Y(n800) );
  MX2 U835 ( .A(\fifo_write/mem[28][3] ), .B(\fifo_write/mem[29][3] ), .S0(
        n1362), .Y(n801) );
  MX2 U836 ( .A(\fifo_write/mem[30][3] ), .B(\fifo_write/mem[31][3] ), .S0(
        n1363), .Y(n802) );
  MX2 U837 ( .A(n787), .B(n788), .S0(n1184), .Y(n803) );
  MX2 U838 ( .A(n789), .B(n790), .S0(n1341), .Y(n804) );
  MX2 U839 ( .A(n791), .B(n792), .S0(n1341), .Y(n805) );
  MX2 U840 ( .A(n793), .B(n794), .S0(n1341), .Y(n806) );
  MX2 U841 ( .A(n795), .B(n796), .S0(n1183), .Y(n807) );
  MX2 U842 ( .A(n797), .B(n798), .S0(\fifo_write/rbin[1] ), .Y(n808) );
  MX2 U843 ( .A(n799), .B(n800), .S0(n1184), .Y(n809) );
  MX2 U844 ( .A(n801), .B(n802), .S0(n1183), .Y(n810) );
  MX2 U845 ( .A(n803), .B(n804), .S0(n1347), .Y(n811) );
  MX2 U846 ( .A(n805), .B(n806), .S0(\fifo_write/rbin[2] ), .Y(n812) );
  MX2 U847 ( .A(n807), .B(n808), .S0(n1348), .Y(n813) );
  MX2 U848 ( .A(n809), .B(n810), .S0(n1347), .Y(n814) );
  MX2 U849 ( .A(n811), .B(n812), .S0(n1332), .Y(n815) );
  MX2 U850 ( .A(n813), .B(n814), .S0(n1332), .Y(n816) );
  MX2 U851 ( .A(n815), .B(n816), .S0(n1188), .Y(wdata_to_fifo[3]) );
  MX2 U852 ( .A(\fifo_write/mem[0][4] ), .B(\fifo_write/mem[1][4] ), .S0(n1363), .Y(n817) );
  MX2 U853 ( .A(\fifo_write/mem[2][4] ), .B(\fifo_write/mem[3][4] ), .S0(n1363), .Y(n818) );
  MX2 U854 ( .A(\fifo_write/mem[4][4] ), .B(\fifo_write/mem[5][4] ), .S0(n1363), .Y(n819) );
  MX2 U855 ( .A(\fifo_write/mem[6][4] ), .B(\fifo_write/mem[7][4] ), .S0(n1363), .Y(n820) );
  MX2 U856 ( .A(\fifo_write/mem[8][4] ), .B(\fifo_write/mem[9][4] ), .S0(n1363), .Y(n821) );
  MX2 U857 ( .A(\fifo_write/mem[10][4] ), .B(\fifo_write/mem[11][4] ), .S0(
        n1363), .Y(n822) );
  MX2 U858 ( .A(\fifo_write/mem[12][4] ), .B(\fifo_write/mem[13][4] ), .S0(
        n1363), .Y(n823) );
  MX2 U859 ( .A(\fifo_write/mem[14][4] ), .B(\fifo_write/mem[15][4] ), .S0(
        n1363), .Y(n824) );
  MX2 U860 ( .A(\fifo_write/mem[16][4] ), .B(\fifo_write/mem[17][4] ), .S0(
        n1364), .Y(n825) );
  MX2 U861 ( .A(\fifo_write/mem[18][4] ), .B(\fifo_write/mem[19][4] ), .S0(
        n1364), .Y(n826) );
  MX2 U862 ( .A(\fifo_write/mem[20][4] ), .B(\fifo_write/mem[21][4] ), .S0(
        n1364), .Y(n827) );
  MX2 U863 ( .A(\fifo_write/mem[22][4] ), .B(\fifo_write/mem[23][4] ), .S0(
        n1364), .Y(n828) );
  MX2 U864 ( .A(\fifo_write/mem[24][4] ), .B(\fifo_write/mem[25][4] ), .S0(
        n1364), .Y(n829) );
  MX2 U865 ( .A(\fifo_write/mem[26][4] ), .B(\fifo_write/mem[27][4] ), .S0(
        n1364), .Y(n830) );
  MX2 U866 ( .A(\fifo_write/mem[28][4] ), .B(\fifo_write/mem[29][4] ), .S0(
        n1364), .Y(n831) );
  MX2 U867 ( .A(\fifo_write/mem[30][4] ), .B(\fifo_write/mem[31][4] ), .S0(
        n1364), .Y(n832) );
  MX2 U868 ( .A(n817), .B(n818), .S0(n1184), .Y(n833) );
  MX2 U869 ( .A(n819), .B(n820), .S0(n1184), .Y(n834) );
  MX2 U870 ( .A(n821), .B(n822), .S0(n1184), .Y(n835) );
  MX2 U871 ( .A(n823), .B(n824), .S0(n1183), .Y(n836) );
  MX2 U872 ( .A(n825), .B(n826), .S0(n1183), .Y(n837) );
  MX2 U873 ( .A(n827), .B(n828), .S0(n1342), .Y(n838) );
  MX2 U874 ( .A(n829), .B(n830), .S0(n1342), .Y(n839) );
  MX2 U875 ( .A(n831), .B(n832), .S0(n1342), .Y(n840) );
  MX2 U876 ( .A(n833), .B(n834), .S0(\fifo_write/rbin[2] ), .Y(n841) );
  MX2 U877 ( .A(n835), .B(n836), .S0(n1348), .Y(n842) );
  MX2 U878 ( .A(n837), .B(n838), .S0(n1347), .Y(n843) );
  MX2 U879 ( .A(n839), .B(n840), .S0(n1348), .Y(n844) );
  MX2 U880 ( .A(n841), .B(n842), .S0(n1332), .Y(n845) );
  MX2 U881 ( .A(n843), .B(n844), .S0(n1332), .Y(n846) );
  MX2 U882 ( .A(n845), .B(n846), .S0(n1188), .Y(wdata_to_fifo[4]) );
  MX2 U883 ( .A(\fifo_write/mem[0][5] ), .B(\fifo_write/mem[1][5] ), .S0(n1364), .Y(n847) );
  MX2 U884 ( .A(\fifo_write/mem[2][5] ), .B(\fifo_write/mem[3][5] ), .S0(n1365), .Y(n848) );
  MX2 U885 ( .A(\fifo_write/mem[4][5] ), .B(\fifo_write/mem[5][5] ), .S0(n1365), .Y(n849) );
  MX2 U886 ( .A(\fifo_write/mem[6][5] ), .B(\fifo_write/mem[7][5] ), .S0(n1365), .Y(n850) );
  MX2 U887 ( .A(\fifo_write/mem[8][5] ), .B(\fifo_write/mem[9][5] ), .S0(n1365), .Y(n851) );
  MX2 U888 ( .A(\fifo_write/mem[10][5] ), .B(\fifo_write/mem[11][5] ), .S0(
        n1365), .Y(n852) );
  MX2 U889 ( .A(\fifo_write/mem[12][5] ), .B(\fifo_write/mem[13][5] ), .S0(
        n1365), .Y(n853) );
  MX2 U890 ( .A(\fifo_write/mem[14][5] ), .B(\fifo_write/mem[15][5] ), .S0(
        n1365), .Y(n854) );
  MX2 U891 ( .A(\fifo_write/mem[16][5] ), .B(\fifo_write/mem[17][5] ), .S0(
        n1365), .Y(n855) );
  MX2 U892 ( .A(\fifo_write/mem[18][5] ), .B(\fifo_write/mem[19][5] ), .S0(
        n1365), .Y(n856) );
  MX2 U893 ( .A(\fifo_write/mem[20][5] ), .B(\fifo_write/mem[21][5] ), .S0(
        n1366), .Y(n857) );
  MX2 U894 ( .A(\fifo_write/mem[22][5] ), .B(\fifo_write/mem[23][5] ), .S0(
        n1366), .Y(n858) );
  MX2 U895 ( .A(\fifo_write/mem[24][5] ), .B(\fifo_write/mem[25][5] ), .S0(
        n1366), .Y(n859) );
  MX2 U896 ( .A(\fifo_write/mem[26][5] ), .B(\fifo_write/mem[27][5] ), .S0(
        n1366), .Y(n860) );
  MX2 U897 ( .A(\fifo_write/mem[28][5] ), .B(\fifo_write/mem[29][5] ), .S0(
        n1366), .Y(n861) );
  MX2 U898 ( .A(\fifo_write/mem[30][5] ), .B(\fifo_write/mem[31][5] ), .S0(
        n1366), .Y(n862) );
  MX2 U899 ( .A(n847), .B(n848), .S0(n1184), .Y(n863) );
  MX2 U900 ( .A(n849), .B(n850), .S0(n1341), .Y(n864) );
  MX2 U901 ( .A(n851), .B(n852), .S0(n1341), .Y(n865) );
  MX2 U902 ( .A(n853), .B(n854), .S0(n1341), .Y(n866) );
  MX2 U903 ( .A(n855), .B(n856), .S0(n1183), .Y(n867) );
  MX2 U904 ( .A(n857), .B(n858), .S0(\fifo_write/rbin[1] ), .Y(n868) );
  MX2 U905 ( .A(n859), .B(n860), .S0(\fifo_write/rbin[1] ), .Y(n869) );
  MX2 U906 ( .A(n861), .B(n862), .S0(n1184), .Y(n870) );
  MX2 U907 ( .A(n863), .B(n864), .S0(n1348), .Y(n871) );
  MX2 U908 ( .A(n865), .B(n866), .S0(n1347), .Y(n872) );
  MX2 U909 ( .A(n867), .B(n868), .S0(n1347), .Y(n873) );
  MX2 U910 ( .A(n869), .B(n870), .S0(n1348), .Y(n874) );
  MX2 U911 ( .A(n871), .B(n872), .S0(n1332), .Y(n875) );
  MX2 U912 ( .A(n873), .B(n874), .S0(n1332), .Y(n876) );
  MX2 U913 ( .A(n875), .B(n876), .S0(n1188), .Y(wdata_to_fifo[5]) );
  MX2 U914 ( .A(\fifo_write/mem[0][6] ), .B(\fifo_write/mem[1][6] ), .S0(n1366), .Y(n877) );
  MX2 U915 ( .A(\fifo_write/mem[2][6] ), .B(\fifo_write/mem[3][6] ), .S0(n1366), .Y(n878) );
  MX2 U916 ( .A(\fifo_write/mem[4][6] ), .B(\fifo_write/mem[5][6] ), .S0(n1366), .Y(n879) );
  MX2 U917 ( .A(\fifo_write/mem[6][6] ), .B(\fifo_write/mem[7][6] ), .S0(n1364), .Y(n880) );
  MX2 U918 ( .A(\fifo_write/mem[8][6] ), .B(\fifo_write/mem[9][6] ), .S0(n1362), .Y(n881) );
  MX2 U919 ( .A(\fifo_write/mem[10][6] ), .B(\fifo_write/mem[11][6] ), .S0(
        n1359), .Y(n882) );
  MX2 U920 ( .A(\fifo_write/mem[12][6] ), .B(\fifo_write/mem[13][6] ), .S0(
        n1361), .Y(n883) );
  MX2 U921 ( .A(\fifo_write/mem[14][6] ), .B(\fifo_write/mem[15][6] ), .S0(
        n1367), .Y(n884) );
  MX2 U922 ( .A(\fifo_write/mem[16][6] ), .B(\fifo_write/mem[17][6] ), .S0(
        n1363), .Y(n885) );
  MX2 U923 ( .A(\fifo_write/mem[18][6] ), .B(\fifo_write/mem[19][6] ), .S0(
        n1360), .Y(n886) );
  MX2 U924 ( .A(\fifo_write/mem[20][6] ), .B(\fifo_write/mem[21][6] ), .S0(
        n1366), .Y(n887) );
  MX2 U925 ( .A(\fifo_write/mem[22][6] ), .B(\fifo_write/mem[23][6] ), .S0(
        n1365), .Y(n888) );
  MX2 U926 ( .A(\fifo_write/mem[24][6] ), .B(\fifo_write/mem[25][6] ), .S0(
        n1361), .Y(n889) );
  MX2 U927 ( .A(\fifo_write/mem[26][6] ), .B(\fifo_write/mem[27][6] ), .S0(
        n1367), .Y(n890) );
  MX2 U928 ( .A(\fifo_write/mem[28][6] ), .B(\fifo_write/mem[29][6] ), .S0(
        n1363), .Y(n891) );
  MX2 U929 ( .A(\fifo_write/mem[30][6] ), .B(\fifo_write/mem[31][6] ), .S0(
        n1360), .Y(n892) );
  MX2 U930 ( .A(n877), .B(n878), .S0(n1184), .Y(n893) );
  MX2 U931 ( .A(n879), .B(n880), .S0(n1183), .Y(n894) );
  MX2 U932 ( .A(n881), .B(n882), .S0(n1341), .Y(n895) );
  MX2 U933 ( .A(n883), .B(n884), .S0(n1342), .Y(n896) );
  MX2 U934 ( .A(n885), .B(n886), .S0(n1183), .Y(n897) );
  MX2 U935 ( .A(n887), .B(n888), .S0(n1342), .Y(n898) );
  MX2 U936 ( .A(n889), .B(n890), .S0(n1342), .Y(n899) );
  MX2 U937 ( .A(n891), .B(n892), .S0(n1342), .Y(n900) );
  MX2 U938 ( .A(n893), .B(n894), .S0(n1347), .Y(n901) );
  MX2 U939 ( .A(n895), .B(n896), .S0(n1348), .Y(n902) );
  MX2 U940 ( .A(n897), .B(n898), .S0(n1348), .Y(n903) );
  MX2 U941 ( .A(n899), .B(n900), .S0(n1347), .Y(n904) );
  MX2 U942 ( .A(n901), .B(n902), .S0(\fifo_write/rbin[3] ), .Y(n905) );
  MX2 U943 ( .A(n903), .B(n904), .S0(n1332), .Y(n906) );
  MX2 U944 ( .A(n905), .B(n906), .S0(n1188), .Y(wdata_to_fifo[6]) );
  MX2 U945 ( .A(\fifo_write/mem[0][7] ), .B(\fifo_write/mem[1][7] ), .S0(n1364), .Y(n907) );
  MX2 U946 ( .A(\fifo_write/mem[2][7] ), .B(\fifo_write/mem[3][7] ), .S0(n1366), .Y(n908) );
  MX2 U947 ( .A(\fifo_write/mem[4][7] ), .B(\fifo_write/mem[5][7] ), .S0(n1365), .Y(n909) );
  MX2 U948 ( .A(\fifo_write/mem[6][7] ), .B(\fifo_write/mem[7][7] ), .S0(n1364), .Y(n910) );
  MX2 U949 ( .A(\fifo_write/mem[8][7] ), .B(\fifo_write/mem[9][7] ), .S0(n1362), .Y(n911) );
  MX2 U950 ( .A(\fifo_write/mem[10][7] ), .B(\fifo_write/mem[11][7] ), .S0(
        n1367), .Y(n912) );
  MX2 U951 ( .A(\fifo_write/mem[12][7] ), .B(\fifo_write/mem[13][7] ), .S0(
        n1363), .Y(n913) );
  MX2 U952 ( .A(\fifo_write/mem[14][7] ), .B(\fifo_write/mem[15][7] ), .S0(
        n1360), .Y(n914) );
  MX2 U953 ( .A(\fifo_write/mem[16][7] ), .B(\fifo_write/mem[17][7] ), .S0(
        n1359), .Y(n915) );
  MX2 U954 ( .A(\fifo_write/mem[18][7] ), .B(\fifo_write/mem[19][7] ), .S0(
        n1362), .Y(n916) );
  MX2 U955 ( .A(\fifo_write/mem[20][7] ), .B(\fifo_write/mem[21][7] ), .S0(
        n1366), .Y(n917) );
  MX2 U956 ( .A(\fifo_write/mem[22][7] ), .B(\fifo_write/mem[23][7] ), .S0(
        n1365), .Y(n918) );
  MX2 U957 ( .A(\fifo_write/mem[24][7] ), .B(\fifo_write/mem[25][7] ), .S0(
        n1364), .Y(n919) );
  MX2 U958 ( .A(\fifo_write/mem[26][7] ), .B(\fifo_write/mem[27][7] ), .S0(
        n1362), .Y(n920) );
  MX2 U959 ( .A(\fifo_write/mem[28][7] ), .B(\fifo_write/mem[29][7] ), .S0(
        n1367), .Y(n921) );
  MX2 U960 ( .A(\fifo_write/mem[30][7] ), .B(\fifo_write/mem[31][7] ), .S0(
        n1367), .Y(n922) );
  MX2 U961 ( .A(n907), .B(n908), .S0(n1184), .Y(n923) );
  MX2 U962 ( .A(n909), .B(n910), .S0(n1341), .Y(n924) );
  MX2 U963 ( .A(n911), .B(n912), .S0(n1341), .Y(n925) );
  MX2 U964 ( .A(n913), .B(n914), .S0(n1341), .Y(n926) );
  MX2 U965 ( .A(n915), .B(n916), .S0(n1183), .Y(n927) );
  MX2 U966 ( .A(n917), .B(n918), .S0(\fifo_write/rbin[1] ), .Y(n928) );
  MX2 U967 ( .A(n919), .B(n920), .S0(\fifo_write/rbin[1] ), .Y(n929) );
  MX2 U968 ( .A(n921), .B(n922), .S0(n1183), .Y(n930) );
  MX2 U969 ( .A(n923), .B(n924), .S0(n1347), .Y(n931) );
  MX2 U970 ( .A(n925), .B(n926), .S0(n1348), .Y(n932) );
  MX2 U971 ( .A(n927), .B(n928), .S0(n1347), .Y(n933) );
  MX2 U972 ( .A(n929), .B(n930), .S0(n1348), .Y(n934) );
  MX2 U973 ( .A(n931), .B(n932), .S0(\fifo_write/rbin[3] ), .Y(n935) );
  MX2 U974 ( .A(n933), .B(n934), .S0(n1332), .Y(n936) );
  MX2 U975 ( .A(n935), .B(n936), .S0(n1188), .Y(wdata_to_fifo[7]) );
  MX2 U976 ( .A(\fifo_read/mem[0][0] ), .B(\fifo_read/mem[1][0] ), .S0(n1351), 
        .Y(n937) );
  MX2 U977 ( .A(\fifo_read/mem[2][0] ), .B(\fifo_read/mem[3][0] ), .S0(n1357), 
        .Y(n938) );
  MX2 U978 ( .A(\fifo_read/mem[4][0] ), .B(\fifo_read/mem[5][0] ), .S0(n1353), 
        .Y(n939) );
  MX2 U979 ( .A(\fifo_read/mem[6][0] ), .B(\fifo_read/mem[7][0] ), .S0(n1349), 
        .Y(n940) );
  MX2 U980 ( .A(\fifo_read/mem[8][0] ), .B(\fifo_read/mem[9][0] ), .S0(n1351), 
        .Y(n941) );
  MX2 U981 ( .A(\fifo_read/mem[10][0] ), .B(\fifo_read/mem[11][0] ), .S0(n1349), .Y(n942) );
  MX2 U982 ( .A(\fifo_read/mem[12][0] ), .B(\fifo_read/mem[13][0] ), .S0(n1356), .Y(n943) );
  MX2 U983 ( .A(\fifo_read/mem[14][0] ), .B(\fifo_read/mem[15][0] ), .S0(n1355), .Y(n944) );
  MX2 U984 ( .A(\fifo_read/mem[16][0] ), .B(\fifo_read/mem[17][0] ), .S0(n1354), .Y(n945) );
  MX2 U985 ( .A(\fifo_read/mem[18][0] ), .B(\fifo_read/mem[19][0] ), .S0(n1352), .Y(n946) );
  MX2 U986 ( .A(\fifo_read/mem[20][0] ), .B(\fifo_read/mem[21][0] ), .S0(n1349), .Y(n947) );
  MX2 U987 ( .A(\fifo_read/mem[22][0] ), .B(\fifo_read/mem[23][0] ), .S0(n1350), .Y(n948) );
  MX2 U988 ( .A(\fifo_read/mem[24][0] ), .B(\fifo_read/mem[25][0] ), .S0(n1351), .Y(n949) );
  MX2 U989 ( .A(\fifo_read/mem[26][0] ), .B(\fifo_read/mem[27][0] ), .S0(n1357), .Y(n950) );
  MX2 U990 ( .A(\fifo_read/mem[28][0] ), .B(\fifo_read/mem[29][0] ), .S0(n1357), .Y(n951) );
  MX2 U991 ( .A(\fifo_read/mem[30][0] ), .B(\fifo_read/mem[31][0] ), .S0(n1357), .Y(n952) );
  MX2 U992 ( .A(n937), .B(n938), .S0(n1182), .Y(n953) );
  MX2 U993 ( .A(n939), .B(n940), .S0(n1339), .Y(n954) );
  MX2 U994 ( .A(n941), .B(n942), .S0(n1339), .Y(n955) );
  MX2 U995 ( .A(n943), .B(n944), .S0(n1338), .Y(n956) );
  MX2 U996 ( .A(n945), .B(n946), .S0(n1181), .Y(n957) );
  MX2 U997 ( .A(n947), .B(n948), .S0(n1339), .Y(n958) );
  MX2 U998 ( .A(n949), .B(n950), .S0(n1339), .Y(n959) );
  MX2 U999 ( .A(n951), .B(n952), .S0(n1339), .Y(n960) );
  MX2 U1000 ( .A(n953), .B(n954), .S0(n1344), .Y(n961) );
  MX2 U1001 ( .A(n955), .B(n956), .S0(\fifo_read/rbin[2] ), .Y(n962) );
  MX2 U1002 ( .A(n957), .B(n958), .S0(n1345), .Y(n963) );
  MX2 U1003 ( .A(n959), .B(n960), .S0(n1344), .Y(n964) );
  MX2 U1004 ( .A(n961), .B(n962), .S0(\fifo_read/rbin[3] ), .Y(n965) );
  MX2 U1005 ( .A(n963), .B(n964), .S0(n1330), .Y(n966) );
  MX2 U1006 ( .A(n965), .B(n966), .S0(n1186), .Y(o_rdata[0]) );
  MX2 U1007 ( .A(\fifo_read/mem[0][1] ), .B(\fifo_read/mem[1][1] ), .S0(n1357), 
        .Y(n967) );
  MX2 U1008 ( .A(\fifo_read/mem[2][1] ), .B(\fifo_read/mem[3][1] ), .S0(
        \fifo_read/rbin[0] ), .Y(n968) );
  MX2 U1009 ( .A(\fifo_read/mem[4][1] ), .B(\fifo_read/mem[5][1] ), .S0(n1357), 
        .Y(n969) );
  MX2 U1010 ( .A(\fifo_read/mem[6][1] ), .B(\fifo_read/mem[7][1] ), .S0(
        \fifo_read/rbin[0] ), .Y(n970) );
  MX2 U1011 ( .A(\fifo_read/mem[8][1] ), .B(\fifo_read/mem[9][1] ), .S0(n1357), 
        .Y(n971) );
  MX2 U1012 ( .A(\fifo_read/mem[10][1] ), .B(\fifo_read/mem[11][1] ), .S0(
        \fifo_read/rbin[0] ), .Y(n972) );
  MX2 U1013 ( .A(\fifo_read/mem[12][1] ), .B(\fifo_read/mem[13][1] ), .S0(
        n1357), .Y(n973) );
  MX2 U1014 ( .A(\fifo_read/mem[14][1] ), .B(\fifo_read/mem[15][1] ), .S0(
        \fifo_read/rbin[0] ), .Y(n974) );
  MX2 U1015 ( .A(\fifo_read/mem[16][1] ), .B(\fifo_read/mem[17][1] ), .S0(
        n1357), .Y(n975) );
  MX2 U1016 ( .A(\fifo_read/mem[18][1] ), .B(\fifo_read/mem[19][1] ), .S0(
        \fifo_read/rbin[0] ), .Y(n976) );
  MX2 U1017 ( .A(\fifo_read/mem[20][1] ), .B(\fifo_read/mem[21][1] ), .S0(
        \fifo_read/rbin[0] ), .Y(n977) );
  MX2 U1018 ( .A(\fifo_read/mem[22][1] ), .B(\fifo_read/mem[23][1] ), .S0(
        n1349), .Y(n978) );
  MX2 U1019 ( .A(\fifo_read/mem[24][1] ), .B(\fifo_read/mem[25][1] ), .S0(
        n1349), .Y(n979) );
  MX2 U1020 ( .A(\fifo_read/mem[26][1] ), .B(\fifo_read/mem[27][1] ), .S0(
        n1349), .Y(n980) );
  MX2 U1021 ( .A(\fifo_read/mem[28][1] ), .B(\fifo_read/mem[29][1] ), .S0(
        n1349), .Y(n981) );
  MX2 U1022 ( .A(\fifo_read/mem[30][1] ), .B(\fifo_read/mem[31][1] ), .S0(
        n1349), .Y(n982) );
  MX2 U1023 ( .A(n967), .B(n968), .S0(n1182), .Y(n983) );
  MX2 U1024 ( .A(n969), .B(n970), .S0(n1338), .Y(n984) );
  MX2 U1025 ( .A(n971), .B(n972), .S0(n1338), .Y(n985) );
  MX2 U1026 ( .A(n973), .B(n974), .S0(n1338), .Y(n986) );
  MX2 U1027 ( .A(n975), .B(n976), .S0(n1181), .Y(n987) );
  MX2 U1028 ( .A(n977), .B(n978), .S0(\fifo_read/rbin[1] ), .Y(n988) );
  MX2 U1029 ( .A(n979), .B(n980), .S0(n1182), .Y(n989) );
  MX2 U1030 ( .A(n981), .B(n982), .S0(n1182), .Y(n990) );
  MX2 U1031 ( .A(n983), .B(n984), .S0(\fifo_read/rbin[2] ), .Y(n991) );
  MX2 U1032 ( .A(n985), .B(n986), .S0(n1345), .Y(n992) );
  MX2 U1033 ( .A(n987), .B(n988), .S0(n1344), .Y(n993) );
  MX2 U1034 ( .A(n989), .B(n990), .S0(\fifo_read/rbin[2] ), .Y(n994) );
  MX2 U1035 ( .A(n991), .B(n992), .S0(n1330), .Y(n995) );
  MX2 U1036 ( .A(n993), .B(n994), .S0(n1330), .Y(n996) );
  MX2 U1037 ( .A(n995), .B(n996), .S0(n1186), .Y(o_rdata[1]) );
  MX2 U1038 ( .A(\fifo_read/mem[0][2] ), .B(\fifo_read/mem[1][2] ), .S0(n1349), 
        .Y(n997) );
  MX2 U1039 ( .A(\fifo_read/mem[2][2] ), .B(\fifo_read/mem[3][2] ), .S0(n1349), 
        .Y(n998) );
  MX2 U1040 ( .A(\fifo_read/mem[4][2] ), .B(\fifo_read/mem[5][2] ), .S0(n1349), 
        .Y(n999) );
  MX2 U1041 ( .A(\fifo_read/mem[6][2] ), .B(\fifo_read/mem[7][2] ), .S0(n1349), 
        .Y(n1000) );
  MX2 U1042 ( .A(\fifo_read/mem[8][2] ), .B(\fifo_read/mem[9][2] ), .S0(n1350), 
        .Y(n1001) );
  MX2 U1043 ( .A(\fifo_read/mem[10][2] ), .B(\fifo_read/mem[11][2] ), .S0(
        n1350), .Y(n1002) );
  MX2 U1044 ( .A(\fifo_read/mem[12][2] ), .B(\fifo_read/mem[13][2] ), .S0(
        n1350), .Y(n1003) );
  MX2 U1045 ( .A(\fifo_read/mem[14][2] ), .B(\fifo_read/mem[15][2] ), .S0(
        n1350), .Y(n1004) );
  MX2 U1046 ( .A(\fifo_read/mem[16][2] ), .B(\fifo_read/mem[17][2] ), .S0(
        n1350), .Y(n1005) );
  MX2 U1047 ( .A(\fifo_read/mem[18][2] ), .B(\fifo_read/mem[19][2] ), .S0(
        n1350), .Y(n1006) );
  MX2 U1048 ( .A(\fifo_read/mem[20][2] ), .B(\fifo_read/mem[21][2] ), .S0(
        n1350), .Y(n1007) );
  MX2 U1049 ( .A(\fifo_read/mem[22][2] ), .B(\fifo_read/mem[23][2] ), .S0(
        n1350), .Y(n1008) );
  MX2 U1050 ( .A(\fifo_read/mem[24][2] ), .B(\fifo_read/mem[25][2] ), .S0(
        n1350), .Y(n1009) );
  MX2 U1051 ( .A(\fifo_read/mem[26][2] ), .B(\fifo_read/mem[27][2] ), .S0(
        n1351), .Y(n1010) );
  MX2 U1052 ( .A(\fifo_read/mem[28][2] ), .B(\fifo_read/mem[29][2] ), .S0(
        n1351), .Y(n1011) );
  MX2 U1053 ( .A(\fifo_read/mem[30][2] ), .B(\fifo_read/mem[31][2] ), .S0(
        n1351), .Y(n1012) );
  MX2 U1054 ( .A(n997), .B(n998), .S0(n1182), .Y(n1013) );
  MX2 U1055 ( .A(n999), .B(n1000), .S0(n1181), .Y(n1014) );
  MX2 U1056 ( .A(n1001), .B(n1002), .S0(n1181), .Y(n1015) );
  MX2 U1057 ( .A(n1003), .B(n1004), .S0(n1182), .Y(n1016) );
  MX2 U1058 ( .A(n1005), .B(n1006), .S0(n1181), .Y(n1017) );
  MX2 U1059 ( .A(n1007), .B(n1008), .S0(n1339), .Y(n1018) );
  MX2 U1060 ( .A(n1009), .B(n1010), .S0(n1339), .Y(n1019) );
  MX2 U1061 ( .A(n1011), .B(n1012), .S0(n1339), .Y(n1020) );
  MX2 U1062 ( .A(n1013), .B(n1014), .S0(n1345), .Y(n1021) );
  MX2 U1063 ( .A(n1015), .B(n1016), .S0(n1344), .Y(n1022) );
  MX2 U1064 ( .A(n1017), .B(n1018), .S0(\fifo_read/rbin[2] ), .Y(n1023) );
  MX2 U1065 ( .A(n1019), .B(n1020), .S0(n1345), .Y(n1024) );
  MX2 U1066 ( .A(n1021), .B(n1022), .S0(n1330), .Y(n1025) );
  MX2 U1067 ( .A(n1023), .B(n1024), .S0(n1330), .Y(n1026) );
  MX2 U1068 ( .A(n1025), .B(n1026), .S0(n1186), .Y(o_rdata[2]) );
  MX2 U1069 ( .A(\fifo_read/mem[0][3] ), .B(\fifo_read/mem[1][3] ), .S0(n1351), 
        .Y(n1027) );
  MX2 U1070 ( .A(\fifo_read/mem[2][3] ), .B(\fifo_read/mem[3][3] ), .S0(n1351), 
        .Y(n1028) );
  MX2 U1071 ( .A(\fifo_read/mem[4][3] ), .B(\fifo_read/mem[5][3] ), .S0(n1351), 
        .Y(n1029) );
  MX2 U1072 ( .A(\fifo_read/mem[6][3] ), .B(\fifo_read/mem[7][3] ), .S0(n1351), 
        .Y(n1030) );
  MX2 U1073 ( .A(\fifo_read/mem[8][3] ), .B(\fifo_read/mem[9][3] ), .S0(n1351), 
        .Y(n1031) );
  MX2 U1074 ( .A(\fifo_read/mem[10][3] ), .B(\fifo_read/mem[11][3] ), .S0(
        n1351), .Y(n1032) );
  MX2 U1075 ( .A(\fifo_read/mem[12][3] ), .B(\fifo_read/mem[13][3] ), .S0(
        n1352), .Y(n1033) );
  MX2 U1076 ( .A(\fifo_read/mem[14][3] ), .B(\fifo_read/mem[15][3] ), .S0(
        n1352), .Y(n1034) );
  MX2 U1077 ( .A(\fifo_read/mem[16][3] ), .B(\fifo_read/mem[17][3] ), .S0(
        n1352), .Y(n1035) );
  MX2 U1078 ( .A(\fifo_read/mem[18][3] ), .B(\fifo_read/mem[19][3] ), .S0(
        n1352), .Y(n1036) );
  MX2 U1079 ( .A(\fifo_read/mem[20][3] ), .B(\fifo_read/mem[21][3] ), .S0(
        n1352), .Y(n1037) );
  MX2 U1080 ( .A(\fifo_read/mem[22][3] ), .B(\fifo_read/mem[23][3] ), .S0(
        n1352), .Y(n1038) );
  MX2 U1081 ( .A(\fifo_read/mem[24][3] ), .B(\fifo_read/mem[25][3] ), .S0(
        n1352), .Y(n1039) );
  MX2 U1082 ( .A(\fifo_read/mem[26][3] ), .B(\fifo_read/mem[27][3] ), .S0(
        n1352), .Y(n1040) );
  MX2 U1083 ( .A(\fifo_read/mem[28][3] ), .B(\fifo_read/mem[29][3] ), .S0(
        n1352), .Y(n1041) );
  MX2 U1084 ( .A(\fifo_read/mem[30][3] ), .B(\fifo_read/mem[31][3] ), .S0(
        n1353), .Y(n1042) );
  MX2 U1085 ( .A(n1027), .B(n1028), .S0(n1182), .Y(n1043) );
  MX2 U1086 ( .A(n1029), .B(n1030), .S0(n1338), .Y(n1044) );
  MX2 U1087 ( .A(n1031), .B(n1032), .S0(n1338), .Y(n1045) );
  MX2 U1088 ( .A(n1033), .B(n1034), .S0(n1338), .Y(n1046) );
  MX2 U1089 ( .A(n1035), .B(n1036), .S0(n1181), .Y(n1047) );
  MX2 U1090 ( .A(n1037), .B(n1038), .S0(\fifo_read/rbin[1] ), .Y(n1048) );
  MX2 U1091 ( .A(n1039), .B(n1040), .S0(n1182), .Y(n1049) );
  MX2 U1092 ( .A(n1041), .B(n1042), .S0(n1181), .Y(n1050) );
  MX2 U1093 ( .A(n1043), .B(n1044), .S0(n1344), .Y(n1051) );
  MX2 U1094 ( .A(n1045), .B(n1046), .S0(\fifo_read/rbin[2] ), .Y(n1052) );
  MX2 U1095 ( .A(n1047), .B(n1048), .S0(n1345), .Y(n1053) );
  MX2 U1096 ( .A(n1049), .B(n1050), .S0(n1344), .Y(n1054) );
  MX2 U1097 ( .A(n1051), .B(n1052), .S0(n1330), .Y(n1055) );
  MX2 U1098 ( .A(n1053), .B(n1054), .S0(n1330), .Y(n1056) );
  MX2 U1099 ( .A(n1055), .B(n1056), .S0(n1186), .Y(o_rdata[3]) );
  MX2 U1100 ( .A(\fifo_read/mem[0][4] ), .B(\fifo_read/mem[1][4] ), .S0(n1353), 
        .Y(n1057) );
  MX2 U1101 ( .A(\fifo_read/mem[2][4] ), .B(\fifo_read/mem[3][4] ), .S0(n1353), 
        .Y(n1058) );
  MX2 U1102 ( .A(\fifo_read/mem[4][4] ), .B(\fifo_read/mem[5][4] ), .S0(n1353), 
        .Y(n1059) );
  MX2 U1103 ( .A(\fifo_read/mem[6][4] ), .B(\fifo_read/mem[7][4] ), .S0(n1353), 
        .Y(n1060) );
  MX2 U1104 ( .A(\fifo_read/mem[8][4] ), .B(\fifo_read/mem[9][4] ), .S0(n1353), 
        .Y(n1061) );
  MX2 U1105 ( .A(\fifo_read/mem[10][4] ), .B(\fifo_read/mem[11][4] ), .S0(
        n1353), .Y(n1062) );
  MX2 U1106 ( .A(\fifo_read/mem[12][4] ), .B(\fifo_read/mem[13][4] ), .S0(
        n1353), .Y(n1063) );
  MX2 U1107 ( .A(\fifo_read/mem[14][4] ), .B(\fifo_read/mem[15][4] ), .S0(
        n1353), .Y(n1064) );
  MX2 U1108 ( .A(\fifo_read/mem[16][4] ), .B(\fifo_read/mem[17][4] ), .S0(
        n1354), .Y(n1065) );
  MX2 U1109 ( .A(\fifo_read/mem[18][4] ), .B(\fifo_read/mem[19][4] ), .S0(
        n1354), .Y(n1066) );
  MX2 U1110 ( .A(\fifo_read/mem[20][4] ), .B(\fifo_read/mem[21][4] ), .S0(
        n1354), .Y(n1067) );
  MX2 U1111 ( .A(\fifo_read/mem[22][4] ), .B(\fifo_read/mem[23][4] ), .S0(
        n1354), .Y(n1068) );
  MX2 U1112 ( .A(\fifo_read/mem[24][4] ), .B(\fifo_read/mem[25][4] ), .S0(
        n1354), .Y(n1069) );
  MX2 U1113 ( .A(\fifo_read/mem[26][4] ), .B(\fifo_read/mem[27][4] ), .S0(
        n1354), .Y(n1070) );
  MX2 U1114 ( .A(\fifo_read/mem[28][4] ), .B(\fifo_read/mem[29][4] ), .S0(
        n1354), .Y(n1071) );
  MX2 U1115 ( .A(\fifo_read/mem[30][4] ), .B(\fifo_read/mem[31][4] ), .S0(
        n1354), .Y(n1072) );
  MX2 U1116 ( .A(n1057), .B(n1058), .S0(n1182), .Y(n1073) );
  MX2 U1117 ( .A(n1059), .B(n1060), .S0(n1182), .Y(n1074) );
  MX2 U1118 ( .A(n1061), .B(n1062), .S0(n1182), .Y(n1075) );
  MX2 U1119 ( .A(n1063), .B(n1064), .S0(n1181), .Y(n1076) );
  MX2 U1120 ( .A(n1065), .B(n1066), .S0(n1181), .Y(n1077) );
  MX2 U1121 ( .A(n1067), .B(n1068), .S0(n1339), .Y(n1078) );
  MX2 U1122 ( .A(n1069), .B(n1070), .S0(n1339), .Y(n1079) );
  MX2 U1123 ( .A(n1071), .B(n1072), .S0(n1339), .Y(n1080) );
  MX2 U1124 ( .A(n1073), .B(n1074), .S0(\fifo_read/rbin[2] ), .Y(n1081) );
  MX2 U1125 ( .A(n1075), .B(n1076), .S0(n1345), .Y(n1082) );
  MX2 U1126 ( .A(n1077), .B(n1078), .S0(n1344), .Y(n1083) );
  MX2 U1127 ( .A(n1079), .B(n1080), .S0(n1345), .Y(n1084) );
  MX2 U1128 ( .A(n1081), .B(n1082), .S0(\fifo_read/rbin[3] ), .Y(n1085) );
  MX2 U1129 ( .A(n1083), .B(n1084), .S0(n1330), .Y(n1086) );
  MX2 U1130 ( .A(n1085), .B(n1086), .S0(n1186), .Y(o_rdata[4]) );
  MX2 U1131 ( .A(\fifo_read/mem[0][5] ), .B(\fifo_read/mem[1][5] ), .S0(n1354), 
        .Y(n1087) );
  MX2 U1132 ( .A(\fifo_read/mem[2][5] ), .B(\fifo_read/mem[3][5] ), .S0(n1355), 
        .Y(n1088) );
  MX2 U1133 ( .A(\fifo_read/mem[4][5] ), .B(\fifo_read/mem[5][5] ), .S0(n1355), 
        .Y(n1089) );
  MX2 U1134 ( .A(\fifo_read/mem[6][5] ), .B(\fifo_read/mem[7][5] ), .S0(n1355), 
        .Y(n1090) );
  MX2 U1135 ( .A(\fifo_read/mem[8][5] ), .B(\fifo_read/mem[9][5] ), .S0(n1355), 
        .Y(n1091) );
  MX2 U1136 ( .A(\fifo_read/mem[10][5] ), .B(\fifo_read/mem[11][5] ), .S0(
        n1355), .Y(n1092) );
  MX2 U1137 ( .A(\fifo_read/mem[12][5] ), .B(\fifo_read/mem[13][5] ), .S0(
        n1355), .Y(n1093) );
  MX2 U1138 ( .A(\fifo_read/mem[14][5] ), .B(\fifo_read/mem[15][5] ), .S0(
        n1355), .Y(n1094) );
  MX2 U1139 ( .A(\fifo_read/mem[16][5] ), .B(\fifo_read/mem[17][5] ), .S0(
        n1355), .Y(n1095) );
  MX2 U1140 ( .A(\fifo_read/mem[18][5] ), .B(\fifo_read/mem[19][5] ), .S0(
        n1355), .Y(n1096) );
  MX2 U1141 ( .A(\fifo_read/mem[20][5] ), .B(\fifo_read/mem[21][5] ), .S0(
        n1356), .Y(n1097) );
  MX2 U1142 ( .A(\fifo_read/mem[22][5] ), .B(\fifo_read/mem[23][5] ), .S0(
        n1356), .Y(n1098) );
  MX2 U1143 ( .A(\fifo_read/mem[24][5] ), .B(\fifo_read/mem[25][5] ), .S0(
        n1356), .Y(n1099) );
  MX2 U1144 ( .A(\fifo_read/mem[26][5] ), .B(\fifo_read/mem[27][5] ), .S0(
        n1356), .Y(n1100) );
  MX2 U1145 ( .A(\fifo_read/mem[28][5] ), .B(\fifo_read/mem[29][5] ), .S0(
        n1356), .Y(n1101) );
  MX2 U1146 ( .A(\fifo_read/mem[30][5] ), .B(\fifo_read/mem[31][5] ), .S0(
        n1356), .Y(n1102) );
  MX2 U1147 ( .A(n1087), .B(n1088), .S0(n1182), .Y(n1103) );
  MX2 U1148 ( .A(n1089), .B(n1090), .S0(n1338), .Y(n1104) );
  MX2 U1149 ( .A(n1091), .B(n1092), .S0(n1338), .Y(n1105) );
  MX2 U1150 ( .A(n1093), .B(n1094), .S0(n1338), .Y(n1106) );
  MX2 U1151 ( .A(n1095), .B(n1096), .S0(n1181), .Y(n1107) );
  MX2 U1152 ( .A(n1097), .B(n1098), .S0(\fifo_read/rbin[1] ), .Y(n1108) );
  MX2 U1153 ( .A(n1099), .B(n1100), .S0(\fifo_read/rbin[1] ), .Y(n1109) );
  MX2 U1154 ( .A(n1101), .B(n1102), .S0(n1182), .Y(n1110) );
  MX2 U1155 ( .A(n1103), .B(n1104), .S0(n1345), .Y(n1111) );
  MX2 U1156 ( .A(n1105), .B(n1106), .S0(n1344), .Y(n1112) );
  MX2 U1157 ( .A(n1107), .B(n1108), .S0(n1344), .Y(n1113) );
  MX2 U1158 ( .A(n1109), .B(n1110), .S0(n1345), .Y(n1114) );
  MX2 U1159 ( .A(n1111), .B(n1112), .S0(\fifo_read/rbin[3] ), .Y(n1115) );
  MX2 U1160 ( .A(n1113), .B(n1114), .S0(n1330), .Y(n1116) );
  MX2 U1161 ( .A(n1115), .B(n1116), .S0(n1186), .Y(o_rdata[5]) );
  MX2 U1162 ( .A(\fifo_read/mem[0][6] ), .B(\fifo_read/mem[1][6] ), .S0(n1356), 
        .Y(n1117) );
  MX2 U1163 ( .A(\fifo_read/mem[2][6] ), .B(\fifo_read/mem[3][6] ), .S0(n1356), 
        .Y(n1118) );
  MX2 U1164 ( .A(\fifo_read/mem[4][6] ), .B(\fifo_read/mem[5][6] ), .S0(n1356), 
        .Y(n1119) );
  MX2 U1165 ( .A(\fifo_read/mem[6][6] ), .B(\fifo_read/mem[7][6] ), .S0(n1354), 
        .Y(n1120) );
  MX2 U1166 ( .A(\fifo_read/mem[8][6] ), .B(\fifo_read/mem[9][6] ), .S0(n1352), 
        .Y(n1121) );
  MX2 U1167 ( .A(\fifo_read/mem[10][6] ), .B(\fifo_read/mem[11][6] ), .S0(
        n1349), .Y(n1122) );
  MX2 U1168 ( .A(\fifo_read/mem[12][6] ), .B(\fifo_read/mem[13][6] ), .S0(
        n1351), .Y(n1123) );
  MX2 U1169 ( .A(\fifo_read/mem[14][6] ), .B(\fifo_read/mem[15][6] ), .S0(
        n1357), .Y(n1124) );
  MX2 U1170 ( .A(\fifo_read/mem[16][6] ), .B(\fifo_read/mem[17][6] ), .S0(
        n1353), .Y(n1125) );
  MX2 U1171 ( .A(\fifo_read/mem[18][6] ), .B(\fifo_read/mem[19][6] ), .S0(
        n1350), .Y(n1126) );
  MX2 U1172 ( .A(\fifo_read/mem[20][6] ), .B(\fifo_read/mem[21][6] ), .S0(
        n1356), .Y(n1127) );
  MX2 U1173 ( .A(\fifo_read/mem[22][6] ), .B(\fifo_read/mem[23][6] ), .S0(
        n1355), .Y(n1128) );
  MX2 U1174 ( .A(\fifo_read/mem[24][6] ), .B(\fifo_read/mem[25][6] ), .S0(
        n1351), .Y(n1129) );
  MX2 U1175 ( .A(\fifo_read/mem[26][6] ), .B(\fifo_read/mem[27][6] ), .S0(
        n1357), .Y(n1130) );
  MX2 U1176 ( .A(\fifo_read/mem[28][6] ), .B(\fifo_read/mem[29][6] ), .S0(
        n1353), .Y(n1131) );
  MX2 U1177 ( .A(\fifo_read/mem[30][6] ), .B(\fifo_read/mem[31][6] ), .S0(
        n1350), .Y(n1132) );
  MX2 U1178 ( .A(n1117), .B(n1118), .S0(n1182), .Y(n1133) );
  MX2 U1179 ( .A(n1119), .B(n1120), .S0(n1181), .Y(n1134) );
  MX2 U1180 ( .A(n1121), .B(n1122), .S0(n1338), .Y(n1135) );
  MX2 U1181 ( .A(n1123), .B(n1124), .S0(n1339), .Y(n1136) );
  MX2 U1182 ( .A(n1125), .B(n1126), .S0(n1181), .Y(n1137) );
  MX2 U1183 ( .A(n1127), .B(n1128), .S0(n1339), .Y(n1138) );
  MX2 U1184 ( .A(n1129), .B(n1130), .S0(n1339), .Y(n1139) );
  MX2 U1185 ( .A(n1131), .B(n1132), .S0(n1339), .Y(n1140) );
  MX2 U1186 ( .A(n1133), .B(n1134), .S0(n1344), .Y(n1141) );
  MX2 U1187 ( .A(n1135), .B(n1136), .S0(n1345), .Y(n1142) );
  MX2 U1188 ( .A(n1137), .B(n1138), .S0(n1345), .Y(n1143) );
  MX2 U1189 ( .A(n1139), .B(n1140), .S0(n1344), .Y(n1144) );
  MX2 U1190 ( .A(n1141), .B(n1142), .S0(\fifo_read/rbin[3] ), .Y(n1145) );
  MX2 U1191 ( .A(n1143), .B(n1144), .S0(n1330), .Y(n1146) );
  MX2 U1192 ( .A(n1145), .B(n1146), .S0(n1186), .Y(o_rdata[6]) );
  MX2 U1193 ( .A(\fifo_read/mem[0][7] ), .B(\fifo_read/mem[1][7] ), .S0(n1354), 
        .Y(n1147) );
  MX2 U1194 ( .A(\fifo_read/mem[2][7] ), .B(\fifo_read/mem[3][7] ), .S0(n1356), 
        .Y(n1148) );
  MX2 U1195 ( .A(\fifo_read/mem[4][7] ), .B(\fifo_read/mem[5][7] ), .S0(n1355), 
        .Y(n1149) );
  MX2 U1196 ( .A(\fifo_read/mem[6][7] ), .B(\fifo_read/mem[7][7] ), .S0(n1354), 
        .Y(n1150) );
  MX2 U1197 ( .A(\fifo_read/mem[8][7] ), .B(\fifo_read/mem[9][7] ), .S0(n1352), 
        .Y(n1151) );
  MX2 U1198 ( .A(\fifo_read/mem[10][7] ), .B(\fifo_read/mem[11][7] ), .S0(
        n1357), .Y(n1152) );
  MX2 U1199 ( .A(\fifo_read/mem[12][7] ), .B(\fifo_read/mem[13][7] ), .S0(
        n1353), .Y(n1153) );
  MX2 U1200 ( .A(\fifo_read/mem[14][7] ), .B(\fifo_read/mem[15][7] ), .S0(
        n1350), .Y(n1154) );
  MX2 U1201 ( .A(\fifo_read/mem[16][7] ), .B(\fifo_read/mem[17][7] ), .S0(
        n1349), .Y(n1155) );
  MX2 U1202 ( .A(\fifo_read/mem[18][7] ), .B(\fifo_read/mem[19][7] ), .S0(
        n1352), .Y(n1156) );
  MX2 U1203 ( .A(\fifo_read/mem[20][7] ), .B(\fifo_read/mem[21][7] ), .S0(
        n1356), .Y(n1157) );
  MX2 U1204 ( .A(\fifo_read/mem[22][7] ), .B(\fifo_read/mem[23][7] ), .S0(
        n1355), .Y(n1158) );
  MX2 U1205 ( .A(\fifo_read/mem[24][7] ), .B(\fifo_read/mem[25][7] ), .S0(
        n1354), .Y(n1159) );
  MX2 U1206 ( .A(\fifo_read/mem[26][7] ), .B(\fifo_read/mem[27][7] ), .S0(
        n1352), .Y(n1160) );
  MX2 U1207 ( .A(\fifo_read/mem[28][7] ), .B(\fifo_read/mem[29][7] ), .S0(
        n1357), .Y(n1161) );
  MX2 U1208 ( .A(\fifo_read/mem[30][7] ), .B(\fifo_read/mem[31][7] ), .S0(
        n1357), .Y(n1162) );
  MX2 U1209 ( .A(n1147), .B(n1148), .S0(n1182), .Y(n1163) );
  MX2 U1210 ( .A(n1149), .B(n1150), .S0(n1338), .Y(n1164) );
  MX2 U1211 ( .A(n1151), .B(n1152), .S0(n1338), .Y(n1165) );
  MX2 U1212 ( .A(n1153), .B(n1154), .S0(n1338), .Y(n1166) );
  MX2 U1213 ( .A(n1155), .B(n1156), .S0(n1181), .Y(n1167) );
  MX2 U1214 ( .A(n1157), .B(n1158), .S0(\fifo_read/rbin[1] ), .Y(n1168) );
  MX2 U1215 ( .A(n1159), .B(n1160), .S0(\fifo_read/rbin[1] ), .Y(n1169) );
  MX2 U1216 ( .A(n1161), .B(n1162), .S0(n1181), .Y(n1170) );
  MX2 U1217 ( .A(n1163), .B(n1164), .S0(n1344), .Y(n1171) );
  MX2 U1218 ( .A(n1165), .B(n1166), .S0(n1345), .Y(n1172) );
  MX2 U1219 ( .A(n1167), .B(n1168), .S0(n1344), .Y(n1173) );
  MX2 U1220 ( .A(n1169), .B(n1170), .S0(n1345), .Y(n1174) );
  MX2 U1221 ( .A(n1171), .B(n1172), .S0(\fifo_read/rbin[3] ), .Y(n1175) );
  MX2 U1222 ( .A(n1173), .B(n1174), .S0(n1330), .Y(n1176) );
  MX2 U1223 ( .A(n1175), .B(n1176), .S0(n1186), .Y(o_rdata[7]) );
  INV U1228 ( .A(n1337), .Y(n1181) );
  INV U1229 ( .A(n1337), .Y(n1182) );
  INV U1230 ( .A(n1340), .Y(n1183) );
  INV U1231 ( .A(n1340), .Y(n1184) );
  INV U1232 ( .A(\fifo_read/rbin[4] ), .Y(n1185) );
  INV U1233 ( .A(n1185), .Y(n1186) );
  INV U1234 ( .A(\fifo_write/rbin[4] ), .Y(n1187) );
  INV U1235 ( .A(n1187), .Y(n1188) );
  INV U1236 ( .A(n1452), .Y(n1189) );
  INV U1237 ( .A(n1189), .Y(n1190) );
  INV U1238 ( .A(n1453), .Y(n1191) );
  INV U1239 ( .A(n1191), .Y(n1192) );
  INV U1240 ( .A(n1454), .Y(n1193) );
  INV U1241 ( .A(n1193), .Y(n1194) );
  INV U1242 ( .A(n1458), .Y(n1195) );
  INV U1243 ( .A(n1195), .Y(n1196) );
  INV U1244 ( .A(n1459), .Y(n1197) );
  INV U1245 ( .A(n1197), .Y(n1198) );
  INV U1246 ( .A(n1460), .Y(n1199) );
  INV U1247 ( .A(n1199), .Y(n1200) );
  INV U1248 ( .A(n1461), .Y(n1201) );
  INV U1249 ( .A(n1201), .Y(n1202) );
  INV U1250 ( .A(n1462), .Y(n1203) );
  INV U1251 ( .A(n1203), .Y(n1204) );
  INV U1252 ( .A(n1463), .Y(n1205) );
  INV U1253 ( .A(n1205), .Y(n1206) );
  INV U1254 ( .A(n1465), .Y(n1207) );
  INV U1255 ( .A(n1207), .Y(n1208) );
  INV U1256 ( .A(n1450), .Y(n1209) );
  INV U1257 ( .A(n1209), .Y(n1210) );
  INV U1258 ( .A(n1451), .Y(n1211) );
  INV U1259 ( .A(n1211), .Y(n1212) );
  INV U1260 ( .A(n1448), .Y(n1213) );
  INV U1261 ( .A(n1213), .Y(n1214) );
  INV U1262 ( .A(n1449), .Y(n1215) );
  INV U1263 ( .A(n1215), .Y(n1216) );
  INV U1264 ( .A(n1445), .Y(n1217) );
  INV U1265 ( .A(n1217), .Y(n1218) );
  INV U1266 ( .A(n1447), .Y(n1219) );
  INV U1267 ( .A(n1219), .Y(n1220) );
  INV U1268 ( .A(n1443), .Y(n1221) );
  INV U1269 ( .A(n1221), .Y(n1222) );
  INV U1270 ( .A(n1444), .Y(n1223) );
  INV U1271 ( .A(n1223), .Y(n1224) );
  INV U1272 ( .A(n1441), .Y(n1225) );
  INV U1273 ( .A(n1225), .Y(n1226) );
  INV U1274 ( .A(n1442), .Y(n1227) );
  INV U1275 ( .A(n1227), .Y(n1228) );
  INV U1276 ( .A(n1439), .Y(n1229) );
  INV U1277 ( .A(n1229), .Y(n1230) );
  INV U1278 ( .A(n1440), .Y(n1231) );
  INV U1279 ( .A(n1231), .Y(n1232) );
  INV U1280 ( .A(n1436), .Y(n1233) );
  INV U1281 ( .A(n1233), .Y(n1234) );
  INV U1282 ( .A(n1438), .Y(n1235) );
  INV U1283 ( .A(n1235), .Y(n1236) );
  INV U1284 ( .A(n1431), .Y(n1237) );
  INV U1285 ( .A(n1237), .Y(n1238) );
  INV U1286 ( .A(n1433), .Y(n1239) );
  INV U1287 ( .A(n1239), .Y(n1240) );
  INV U1288 ( .A(n1427), .Y(n1241) );
  INV U1289 ( .A(n1241), .Y(n1242) );
  INV U1290 ( .A(n1429), .Y(n1243) );
  INV U1291 ( .A(n1243), .Y(n1244) );
  INV U1292 ( .A(n1423), .Y(n1245) );
  INV U1293 ( .A(n1245), .Y(n1246) );
  INV U1294 ( .A(n1425), .Y(n1247) );
  INV U1295 ( .A(n1247), .Y(n1248) );
  INV U1296 ( .A(n1418), .Y(n1249) );
  INV U1297 ( .A(n1249), .Y(n1250) );
  INV U1298 ( .A(n1421), .Y(n1251) );
  INV U1299 ( .A(n1251), .Y(n1252) );
  INV U1300 ( .A(n1414), .Y(n1253) );
  INV U1301 ( .A(n1253), .Y(n1254) );
  INV U1302 ( .A(n1416), .Y(n1255) );
  INV U1303 ( .A(n1255), .Y(n1256) );
  INV U1304 ( .A(n1412), .Y(n1257) );
  INV U1305 ( .A(n1257), .Y(n1258) );
  INV U1306 ( .A(n1413), .Y(n1259) );
  INV U1307 ( .A(n1259), .Y(n1260) );
  INV U1308 ( .A(n1410), .Y(n1261) );
  INV U1309 ( .A(n1261), .Y(n1262) );
  INV U1310 ( .A(n1411), .Y(n1263) );
  INV U1311 ( .A(n1263), .Y(n1264) );
  INV U1312 ( .A(n1403), .Y(n1265) );
  INV U1313 ( .A(n1265), .Y(n1266) );
  INV U1314 ( .A(n1404), .Y(n1267) );
  INV U1315 ( .A(n1267), .Y(n1268) );
  INV U1316 ( .A(n1405), .Y(n1269) );
  INV U1317 ( .A(n1269), .Y(n1270) );
  INV U1318 ( .A(n1409), .Y(n1271) );
  INV U1319 ( .A(n1271), .Y(n1272) );
  INV U1320 ( .A(n1399), .Y(n1273) );
  INV U1321 ( .A(n1273), .Y(n1274) );
  INV U1322 ( .A(n1400), .Y(n1275) );
  INV U1323 ( .A(n1275), .Y(n1276) );
  INV U1324 ( .A(n1401), .Y(n1277) );
  INV U1325 ( .A(n1277), .Y(n1278) );
  INV U1326 ( .A(n1402), .Y(n1279) );
  INV U1327 ( .A(n1279), .Y(n1280) );
  INV U1328 ( .A(n1394), .Y(n1281) );
  INV U1329 ( .A(n1281), .Y(n1282) );
  INV U1330 ( .A(n1395), .Y(n1283) );
  INV U1331 ( .A(n1283), .Y(n1284) );
  INV U1332 ( .A(n1396), .Y(n1285) );
  INV U1333 ( .A(n1285), .Y(n1286) );
  INV U1334 ( .A(n1398), .Y(n1287) );
  INV U1335 ( .A(n1287), .Y(n1288) );
  INV U1336 ( .A(n1390), .Y(n1289) );
  INV U1337 ( .A(n1289), .Y(n1290) );
  INV U1338 ( .A(n1391), .Y(n1291) );
  INV U1339 ( .A(n1291), .Y(n1292) );
  INV U1340 ( .A(n1392), .Y(n1293) );
  INV U1341 ( .A(n1293), .Y(n1294) );
  INV U1342 ( .A(n1393), .Y(n1295) );
  INV U1343 ( .A(n1295), .Y(n1296) );
  INV U1344 ( .A(n1382), .Y(n1297) );
  INV U1345 ( .A(n1297), .Y(n1298) );
  INV U1346 ( .A(n1384), .Y(n1299) );
  INV U1347 ( .A(n1299), .Y(n1300) );
  INV U1348 ( .A(n1387), .Y(n1301) );
  INV U1349 ( .A(n1301), .Y(n1302) );
  INV U1350 ( .A(n1389), .Y(n1303) );
  INV U1351 ( .A(n1303), .Y(n1304) );
  INV U1352 ( .A(n1374), .Y(n1305) );
  INV U1353 ( .A(n1305), .Y(n1306) );
  INV U1354 ( .A(n1376), .Y(n1307) );
  INV U1355 ( .A(n1307), .Y(n1308) );
  INV U1356 ( .A(n1378), .Y(n1309) );
  INV U1357 ( .A(n1309), .Y(n1310) );
  INV U1358 ( .A(n1380), .Y(n1311) );
  INV U1359 ( .A(n1311), .Y(n1312) );
  INV U1360 ( .A(wdata_to_fifo[1]), .Y(n1313) );
  INV U1361 ( .A(n1313), .Y(n1314) );
  INV U1362 ( .A(wdata_to_fifo[0]), .Y(n1315) );
  INV U1363 ( .A(n1315), .Y(n1316) );
  INV U1364 ( .A(n1369), .Y(n1317) );
  INV U1365 ( .A(n1317), .Y(n1318) );
  INV U1366 ( .A(n1372), .Y(n1319) );
  INV U1367 ( .A(n1319), .Y(n1320) );
  INV U1368 ( .A(wdata_to_fifo[5]), .Y(n1321) );
  INV U1369 ( .A(n1321), .Y(n1322) );
  INV U1370 ( .A(wdata_to_fifo[4]), .Y(n1323) );
  INV U1371 ( .A(n1323), .Y(n1324) );
  INV U1372 ( .A(wdata_to_fifo[3]), .Y(n1325) );
  INV U1373 ( .A(n1325), .Y(n1326) );
  INV U1374 ( .A(wdata_to_fifo[2]), .Y(n1327) );
  INV U1375 ( .A(n1327), .Y(n1328) );
  INV U1376 ( .A(\fifo_read/rbin[3] ), .Y(n1329) );
  INV U1377 ( .A(n1329), .Y(n1330) );
  INV U1378 ( .A(\fifo_write/rbin[3] ), .Y(n1331) );
  INV U1379 ( .A(n1331), .Y(n1332) );
  INV U1380 ( .A(wdata_to_fifo[7]), .Y(n1333) );
  INV U1381 ( .A(n1333), .Y(n1334) );
  INV U1382 ( .A(wdata_to_fifo[6]), .Y(n1335) );
  INV U1383 ( .A(n1335), .Y(n1336) );
  INV U1384 ( .A(\fifo_read/rbin[1] ), .Y(n1337) );
  INV U1385 ( .A(n1337), .Y(n1338) );
  INV U1386 ( .A(n1337), .Y(n1339) );
  INV U1387 ( .A(\fifo_write/rbin[1] ), .Y(n1340) );
  INV U1388 ( .A(n1340), .Y(n1341) );
  INV U1389 ( .A(n1340), .Y(n1342) );
  INV U1390 ( .A(\fifo_read/rbin[2] ), .Y(n1343) );
  INV U1391 ( .A(n1343), .Y(n1344) );
  INV U1392 ( .A(n1343), .Y(n1345) );
  INV U1393 ( .A(\fifo_write/rbin[2] ), .Y(n1346) );
  INV U1394 ( .A(n1346), .Y(n1347) );
  INV U1395 ( .A(n1346), .Y(n1348) );
  INV U1396 ( .A(n1358), .Y(n1349) );
  INV U1397 ( .A(n1358), .Y(n1350) );
  INV U1398 ( .A(n1358), .Y(n1351) );
  INV U1399 ( .A(n1358), .Y(n1352) );
  INV U1400 ( .A(n1358), .Y(n1353) );
  INV U1401 ( .A(n1358), .Y(n1354) );
  INV U1402 ( .A(n1358), .Y(n1355) );
  INV U1403 ( .A(n1358), .Y(n1356) );
  INV U1404 ( .A(n1358), .Y(n1357) );
  INV U1405 ( .A(\fifo_read/rbin[0] ), .Y(n1358) );
  INV U1406 ( .A(n1368), .Y(n1359) );
  INV U1407 ( .A(n1368), .Y(n1360) );
  INV U1408 ( .A(n1368), .Y(n1361) );
  INV U1409 ( .A(n1368), .Y(n1362) );
  INV U1410 ( .A(n1368), .Y(n1363) );
  INV U1411 ( .A(n1368), .Y(n1364) );
  INV U1412 ( .A(n1368), .Y(n1365) );
  INV U1413 ( .A(n1368), .Y(n1366) );
  INV U1414 ( .A(n1368), .Y(n1367) );
  INV U1415 ( .A(\fifo_write/rbin[0] ), .Y(n1368) );
  MX2 U1416 ( .A(\fifo_write/mem[31][0] ), .B(i_wdata[0]), .S0(n1318), .Y(n696) );
  MX2 U1417 ( .A(\fifo_write/mem[31][1] ), .B(i_wdata[1]), .S0(n1318), .Y(n695) );
  MX2 U1418 ( .A(\fifo_write/mem[31][2] ), .B(i_wdata[2]), .S0(n1318), .Y(n694) );
  MX2 U1419 ( .A(\fifo_write/mem[31][3] ), .B(i_wdata[3]), .S0(n1318), .Y(n693) );
  MX2 U1420 ( .A(\fifo_write/mem[31][4] ), .B(i_wdata[4]), .S0(n1318), .Y(n692) );
  MX2 U1421 ( .A(\fifo_write/mem[31][5] ), .B(i_wdata[5]), .S0(n1318), .Y(n691) );
  MX2 U1422 ( .A(\fifo_write/mem[31][6] ), .B(i_wdata[6]), .S0(n1318), .Y(n690) );
  MX2 U1423 ( .A(\fifo_write/mem[31][7] ), .B(i_wdata[7]), .S0(n1318), .Y(n689) );
  NOR2B U1424 ( .AN(n1370), .B(n1371), .Y(n1369) );
  MX2 U1425 ( .A(\fifo_write/mem[30][0] ), .B(i_wdata[0]), .S0(n1320), .Y(n688) );
  MX2 U1426 ( .A(\fifo_write/mem[30][1] ), .B(i_wdata[1]), .S0(n1320), .Y(n687) );
  MX2 U1427 ( .A(\fifo_write/mem[30][2] ), .B(i_wdata[2]), .S0(n1320), .Y(n686) );
  MX2 U1428 ( .A(\fifo_write/mem[30][3] ), .B(i_wdata[3]), .S0(n1320), .Y(n685) );
  MX2 U1429 ( .A(\fifo_write/mem[30][4] ), .B(i_wdata[4]), .S0(n1320), .Y(n684) );
  MX2 U1430 ( .A(\fifo_write/mem[30][5] ), .B(i_wdata[5]), .S0(n1320), .Y(n683) );
  MX2 U1431 ( .A(\fifo_write/mem[30][6] ), .B(i_wdata[6]), .S0(n1320), .Y(n682) );
  MX2 U1432 ( .A(\fifo_write/mem[30][7] ), .B(i_wdata[7]), .S0(n1320), .Y(n681) );
  NOR2B U1433 ( .AN(n1373), .B(n1371), .Y(n1372) );
  MX2 U1434 ( .A(\fifo_write/mem[29][0] ), .B(i_wdata[0]), .S0(n1306), .Y(n680) );
  MX2 U1435 ( .A(\fifo_write/mem[29][1] ), .B(i_wdata[1]), .S0(n1306), .Y(n679) );
  MX2 U1436 ( .A(\fifo_write/mem[29][2] ), .B(i_wdata[2]), .S0(n1306), .Y(n678) );
  MX2 U1437 ( .A(\fifo_write/mem[29][3] ), .B(i_wdata[3]), .S0(n1306), .Y(n677) );
  MX2 U1438 ( .A(\fifo_write/mem[29][4] ), .B(i_wdata[4]), .S0(n1306), .Y(n676) );
  MX2 U1439 ( .A(\fifo_write/mem[29][5] ), .B(i_wdata[5]), .S0(n1306), .Y(n675) );
  MX2 U1440 ( .A(\fifo_write/mem[29][6] ), .B(i_wdata[6]), .S0(n1306), .Y(n674) );
  MX2 U1441 ( .A(\fifo_write/mem[29][7] ), .B(i_wdata[7]), .S0(n1306), .Y(n673) );
  NOR2B U1442 ( .AN(n1375), .B(n1371), .Y(n1374) );
  MX2 U1443 ( .A(\fifo_write/mem[28][0] ), .B(i_wdata[0]), .S0(n1308), .Y(n672) );
  MX2 U1444 ( .A(\fifo_write/mem[28][1] ), .B(i_wdata[1]), .S0(n1308), .Y(n671) );
  MX2 U1445 ( .A(\fifo_write/mem[28][2] ), .B(i_wdata[2]), .S0(n1308), .Y(n670) );
  MX2 U1446 ( .A(\fifo_write/mem[28][3] ), .B(i_wdata[3]), .S0(n1308), .Y(n669) );
  MX2 U1447 ( .A(\fifo_write/mem[28][4] ), .B(i_wdata[4]), .S0(n1308), .Y(n668) );
  MX2 U1448 ( .A(\fifo_write/mem[28][5] ), .B(i_wdata[5]), .S0(n1308), .Y(n667) );
  MX2 U1449 ( .A(\fifo_write/mem[28][6] ), .B(i_wdata[6]), .S0(n1308), .Y(n666) );
  MX2 U1450 ( .A(\fifo_write/mem[28][7] ), .B(i_wdata[7]), .S0(n1308), .Y(n665) );
  NOR2B U1451 ( .AN(n1377), .B(n1371), .Y(n1376) );
  MX2 U1452 ( .A(\fifo_write/mem[27][0] ), .B(i_wdata[0]), .S0(n1310), .Y(n664) );
  MX2 U1453 ( .A(\fifo_write/mem[27][1] ), .B(i_wdata[1]), .S0(n1310), .Y(n663) );
  MX2 U1454 ( .A(\fifo_write/mem[27][2] ), .B(i_wdata[2]), .S0(n1310), .Y(n662) );
  MX2 U1455 ( .A(\fifo_write/mem[27][3] ), .B(i_wdata[3]), .S0(n1310), .Y(n661) );
  MX2 U1456 ( .A(\fifo_write/mem[27][4] ), .B(i_wdata[4]), .S0(n1310), .Y(n660) );
  MX2 U1457 ( .A(\fifo_write/mem[27][5] ), .B(i_wdata[5]), .S0(n1310), .Y(n659) );
  MX2 U1458 ( .A(\fifo_write/mem[27][6] ), .B(i_wdata[6]), .S0(n1310), .Y(n658) );
  MX2 U1459 ( .A(\fifo_write/mem[27][7] ), .B(i_wdata[7]), .S0(n1310), .Y(n657) );
  NOR2B U1460 ( .AN(n1379), .B(n1371), .Y(n1378) );
  MX2 U1461 ( .A(\fifo_write/mem[26][0] ), .B(i_wdata[0]), .S0(n1312), .Y(n656) );
  MX2 U1462 ( .A(\fifo_write/mem[26][1] ), .B(i_wdata[1]), .S0(n1312), .Y(n655) );
  MX2 U1463 ( .A(\fifo_write/mem[26][2] ), .B(i_wdata[2]), .S0(n1312), .Y(n654) );
  MX2 U1464 ( .A(\fifo_write/mem[26][3] ), .B(i_wdata[3]), .S0(n1312), .Y(n653) );
  MX2 U1465 ( .A(\fifo_write/mem[26][4] ), .B(i_wdata[4]), .S0(n1312), .Y(n652) );
  MX2 U1466 ( .A(\fifo_write/mem[26][5] ), .B(i_wdata[5]), .S0(n1312), .Y(n651) );
  MX2 U1467 ( .A(\fifo_write/mem[26][6] ), .B(i_wdata[6]), .S0(n1312), .Y(n650) );
  MX2 U1468 ( .A(\fifo_write/mem[26][7] ), .B(i_wdata[7]), .S0(n1312), .Y(n649) );
  NOR2B U1469 ( .AN(n1381), .B(n1371), .Y(n1380) );
  MX2 U1470 ( .A(\fifo_write/mem[25][0] ), .B(i_wdata[0]), .S0(n1298), .Y(n648) );
  MX2 U1471 ( .A(\fifo_write/mem[25][1] ), .B(i_wdata[1]), .S0(n1298), .Y(n647) );
  MX2 U1472 ( .A(\fifo_write/mem[25][2] ), .B(i_wdata[2]), .S0(n1298), .Y(n646) );
  MX2 U1473 ( .A(\fifo_write/mem[25][3] ), .B(i_wdata[3]), .S0(n1298), .Y(n645) );
  MX2 U1474 ( .A(\fifo_write/mem[25][4] ), .B(i_wdata[4]), .S0(n1298), .Y(n644) );
  MX2 U1475 ( .A(\fifo_write/mem[25][5] ), .B(i_wdata[5]), .S0(n1298), .Y(n643) );
  MX2 U1476 ( .A(\fifo_write/mem[25][6] ), .B(i_wdata[6]), .S0(n1298), .Y(n642) );
  MX2 U1477 ( .A(\fifo_write/mem[25][7] ), .B(i_wdata[7]), .S0(n1298), .Y(n641) );
  NOR2B U1478 ( .AN(n1383), .B(n1371), .Y(n1382) );
  MX2 U1479 ( .A(\fifo_write/mem[24][0] ), .B(i_wdata[0]), .S0(n1300), .Y(n640) );
  MX2 U1480 ( .A(\fifo_write/mem[24][1] ), .B(i_wdata[1]), .S0(n1300), .Y(n639) );
  MX2 U1481 ( .A(\fifo_write/mem[24][2] ), .B(i_wdata[2]), .S0(n1300), .Y(n638) );
  MX2 U1482 ( .A(\fifo_write/mem[24][3] ), .B(i_wdata[3]), .S0(n1300), .Y(n637) );
  MX2 U1483 ( .A(\fifo_write/mem[24][4] ), .B(i_wdata[4]), .S0(n1300), .Y(n636) );
  MX2 U1484 ( .A(\fifo_write/mem[24][5] ), .B(i_wdata[5]), .S0(n1300), .Y(n635) );
  MX2 U1485 ( .A(\fifo_write/mem[24][6] ), .B(i_wdata[6]), .S0(n1300), .Y(n634) );
  MX2 U1486 ( .A(\fifo_write/mem[24][7] ), .B(i_wdata[7]), .S0(n1300), .Y(n633) );
  NOR2B U1487 ( .AN(n1385), .B(n1371), .Y(n1384) );
  NAND3 U1488 ( .A(n1386), .B(\fifo_write/waddr[4] ), .C(\fifo_write/waddr[3] ), .Y(n1371) );
  MX2 U1489 ( .A(\fifo_write/mem[23][0] ), .B(i_wdata[0]), .S0(n1302), .Y(n632) );
  MX2 U1490 ( .A(\fifo_write/mem[23][1] ), .B(i_wdata[1]), .S0(n1302), .Y(n631) );
  MX2 U1491 ( .A(\fifo_write/mem[23][2] ), .B(i_wdata[2]), .S0(n1302), .Y(n630) );
  MX2 U1492 ( .A(\fifo_write/mem[23][3] ), .B(i_wdata[3]), .S0(n1302), .Y(n629) );
  MX2 U1493 ( .A(\fifo_write/mem[23][4] ), .B(i_wdata[4]), .S0(n1302), .Y(n628) );
  MX2 U1494 ( .A(\fifo_write/mem[23][5] ), .B(i_wdata[5]), .S0(n1302), .Y(n627) );
  MX2 U1495 ( .A(\fifo_write/mem[23][6] ), .B(i_wdata[6]), .S0(n1302), .Y(n626) );
  MX2 U1496 ( .A(\fifo_write/mem[23][7] ), .B(i_wdata[7]), .S0(n1302), .Y(n625) );
  NOR2B U1497 ( .AN(n1370), .B(n1388), .Y(n1387) );
  MX2 U1498 ( .A(\fifo_write/mem[22][0] ), .B(i_wdata[0]), .S0(n1304), .Y(n624) );
  MX2 U1499 ( .A(\fifo_write/mem[22][1] ), .B(i_wdata[1]), .S0(n1304), .Y(n623) );
  MX2 U1500 ( .A(\fifo_write/mem[22][2] ), .B(i_wdata[2]), .S0(n1304), .Y(n622) );
  MX2 U1501 ( .A(\fifo_write/mem[22][3] ), .B(i_wdata[3]), .S0(n1304), .Y(n621) );
  MX2 U1502 ( .A(\fifo_write/mem[22][4] ), .B(i_wdata[4]), .S0(n1304), .Y(n620) );
  MX2 U1503 ( .A(\fifo_write/mem[22][5] ), .B(i_wdata[5]), .S0(n1304), .Y(n619) );
  MX2 U1504 ( .A(\fifo_write/mem[22][6] ), .B(i_wdata[6]), .S0(n1304), .Y(n618) );
  MX2 U1505 ( .A(\fifo_write/mem[22][7] ), .B(i_wdata[7]), .S0(n1304), .Y(n617) );
  NOR2B U1506 ( .AN(n1373), .B(n1388), .Y(n1389) );
  MX2 U1507 ( .A(\fifo_write/mem[21][0] ), .B(i_wdata[0]), .S0(n1290), .Y(n616) );
  MX2 U1508 ( .A(\fifo_write/mem[21][1] ), .B(i_wdata[1]), .S0(n1290), .Y(n615) );
  MX2 U1509 ( .A(\fifo_write/mem[21][2] ), .B(i_wdata[2]), .S0(n1290), .Y(n614) );
  MX2 U1510 ( .A(\fifo_write/mem[21][3] ), .B(i_wdata[3]), .S0(n1290), .Y(n613) );
  MX2 U1511 ( .A(\fifo_write/mem[21][4] ), .B(i_wdata[4]), .S0(n1290), .Y(n612) );
  MX2 U1512 ( .A(\fifo_write/mem[21][5] ), .B(i_wdata[5]), .S0(n1290), .Y(n611) );
  MX2 U1513 ( .A(\fifo_write/mem[21][6] ), .B(i_wdata[6]), .S0(n1290), .Y(n610) );
  MX2 U1514 ( .A(\fifo_write/mem[21][7] ), .B(i_wdata[7]), .S0(n1290), .Y(n609) );
  NOR2B U1515 ( .AN(n1375), .B(n1388), .Y(n1390) );
  MX2 U1516 ( .A(\fifo_write/mem[20][0] ), .B(i_wdata[0]), .S0(n1292), .Y(n608) );
  MX2 U1517 ( .A(\fifo_write/mem[20][1] ), .B(i_wdata[1]), .S0(n1292), .Y(n607) );
  MX2 U1518 ( .A(\fifo_write/mem[20][2] ), .B(i_wdata[2]), .S0(n1292), .Y(n606) );
  MX2 U1519 ( .A(\fifo_write/mem[20][3] ), .B(i_wdata[3]), .S0(n1292), .Y(n605) );
  MX2 U1520 ( .A(\fifo_write/mem[20][4] ), .B(i_wdata[4]), .S0(n1292), .Y(n604) );
  MX2 U1521 ( .A(\fifo_write/mem[20][5] ), .B(i_wdata[5]), .S0(n1292), .Y(n603) );
  MX2 U1522 ( .A(\fifo_write/mem[20][6] ), .B(i_wdata[6]), .S0(n1292), .Y(n602) );
  MX2 U1523 ( .A(\fifo_write/mem[20][7] ), .B(i_wdata[7]), .S0(n1292), .Y(n601) );
  NOR2B U1524 ( .AN(n1377), .B(n1388), .Y(n1391) );
  MX2 U1525 ( .A(\fifo_write/mem[19][0] ), .B(i_wdata[0]), .S0(n1294), .Y(n600) );
  MX2 U1526 ( .A(\fifo_write/mem[19][1] ), .B(i_wdata[1]), .S0(n1294), .Y(n599) );
  MX2 U1527 ( .A(\fifo_write/mem[19][2] ), .B(i_wdata[2]), .S0(n1294), .Y(n598) );
  MX2 U1528 ( .A(\fifo_write/mem[19][3] ), .B(i_wdata[3]), .S0(n1294), .Y(n597) );
  MX2 U1529 ( .A(\fifo_write/mem[19][4] ), .B(i_wdata[4]), .S0(n1294), .Y(n596) );
  MX2 U1530 ( .A(\fifo_write/mem[19][5] ), .B(i_wdata[5]), .S0(n1294), .Y(n595) );
  MX2 U1531 ( .A(\fifo_write/mem[19][6] ), .B(i_wdata[6]), .S0(n1294), .Y(n594) );
  MX2 U1532 ( .A(\fifo_write/mem[19][7] ), .B(i_wdata[7]), .S0(n1294), .Y(n593) );
  NOR2B U1533 ( .AN(n1379), .B(n1388), .Y(n1392) );
  MX2 U1534 ( .A(\fifo_write/mem[18][0] ), .B(i_wdata[0]), .S0(n1296), .Y(n592) );
  MX2 U1535 ( .A(\fifo_write/mem[18][1] ), .B(i_wdata[1]), .S0(n1296), .Y(n591) );
  MX2 U1536 ( .A(\fifo_write/mem[18][2] ), .B(i_wdata[2]), .S0(n1296), .Y(n590) );
  MX2 U1537 ( .A(\fifo_write/mem[18][3] ), .B(i_wdata[3]), .S0(n1296), .Y(n589) );
  MX2 U1538 ( .A(\fifo_write/mem[18][4] ), .B(i_wdata[4]), .S0(n1296), .Y(n588) );
  MX2 U1539 ( .A(\fifo_write/mem[18][5] ), .B(i_wdata[5]), .S0(n1296), .Y(n587) );
  MX2 U1540 ( .A(\fifo_write/mem[18][6] ), .B(i_wdata[6]), .S0(n1296), .Y(n586) );
  MX2 U1541 ( .A(\fifo_write/mem[18][7] ), .B(i_wdata[7]), .S0(n1296), .Y(n585) );
  NOR2B U1542 ( .AN(n1381), .B(n1388), .Y(n1393) );
  MX2 U1543 ( .A(\fifo_write/mem[17][0] ), .B(i_wdata[0]), .S0(n1282), .Y(n584) );
  MX2 U1544 ( .A(\fifo_write/mem[17][1] ), .B(i_wdata[1]), .S0(n1282), .Y(n583) );
  MX2 U1545 ( .A(\fifo_write/mem[17][2] ), .B(i_wdata[2]), .S0(n1282), .Y(n582) );
  MX2 U1546 ( .A(\fifo_write/mem[17][3] ), .B(i_wdata[3]), .S0(n1282), .Y(n581) );
  MX2 U1547 ( .A(\fifo_write/mem[17][4] ), .B(i_wdata[4]), .S0(n1282), .Y(n580) );
  MX2 U1548 ( .A(\fifo_write/mem[17][5] ), .B(i_wdata[5]), .S0(n1282), .Y(n579) );
  MX2 U1549 ( .A(\fifo_write/mem[17][6] ), .B(i_wdata[6]), .S0(n1282), .Y(n578) );
  MX2 U1550 ( .A(\fifo_write/mem[17][7] ), .B(i_wdata[7]), .S0(n1282), .Y(n577) );
  NOR2B U1551 ( .AN(n1383), .B(n1388), .Y(n1394) );
  MX2 U1552 ( .A(\fifo_write/mem[16][0] ), .B(i_wdata[0]), .S0(n1284), .Y(n576) );
  MX2 U1553 ( .A(\fifo_write/mem[16][1] ), .B(i_wdata[1]), .S0(n1284), .Y(n575) );
  MX2 U1554 ( .A(\fifo_write/mem[16][2] ), .B(i_wdata[2]), .S0(n1284), .Y(n574) );
  MX2 U1555 ( .A(\fifo_write/mem[16][3] ), .B(i_wdata[3]), .S0(n1284), .Y(n573) );
  MX2 U1556 ( .A(\fifo_write/mem[16][4] ), .B(i_wdata[4]), .S0(n1284), .Y(n572) );
  MX2 U1557 ( .A(\fifo_write/mem[16][5] ), .B(i_wdata[5]), .S0(n1284), .Y(n571) );
  MX2 U1558 ( .A(\fifo_write/mem[16][6] ), .B(i_wdata[6]), .S0(n1284), .Y(n570) );
  MX2 U1559 ( .A(\fifo_write/mem[16][7] ), .B(i_wdata[7]), .S0(n1284), .Y(n569) );
  NOR2B U1560 ( .AN(n1385), .B(n1388), .Y(n1395) );
  NAND3B U1561 ( .AN(\fifo_write/waddr[3] ), .B(\fifo_write/waddr[4] ), .C(
        n1386), .Y(n1388) );
  MX2 U1562 ( .A(\fifo_write/mem[15][0] ), .B(i_wdata[0]), .S0(n1286), .Y(n568) );
  MX2 U1563 ( .A(\fifo_write/mem[15][1] ), .B(i_wdata[1]), .S0(n1286), .Y(n567) );
  MX2 U1564 ( .A(\fifo_write/mem[15][2] ), .B(i_wdata[2]), .S0(n1286), .Y(n566) );
  MX2 U1565 ( .A(\fifo_write/mem[15][3] ), .B(i_wdata[3]), .S0(n1286), .Y(n565) );
  MX2 U1566 ( .A(\fifo_write/mem[15][4] ), .B(i_wdata[4]), .S0(n1286), .Y(n564) );
  MX2 U1567 ( .A(\fifo_write/mem[15][5] ), .B(i_wdata[5]), .S0(n1286), .Y(n563) );
  MX2 U1568 ( .A(\fifo_write/mem[15][6] ), .B(i_wdata[6]), .S0(n1286), .Y(n562) );
  MX2 U1569 ( .A(\fifo_write/mem[15][7] ), .B(i_wdata[7]), .S0(n1286), .Y(n561) );
  NOR2B U1570 ( .AN(n1370), .B(n1397), .Y(n1396) );
  MX2 U1571 ( .A(\fifo_write/mem[14][0] ), .B(i_wdata[0]), .S0(n1288), .Y(n560) );
  MX2 U1572 ( .A(\fifo_write/mem[14][1] ), .B(i_wdata[1]), .S0(n1288), .Y(n559) );
  MX2 U1573 ( .A(\fifo_write/mem[14][2] ), .B(i_wdata[2]), .S0(n1288), .Y(n558) );
  MX2 U1574 ( .A(\fifo_write/mem[14][3] ), .B(i_wdata[3]), .S0(n1288), .Y(n557) );
  MX2 U1575 ( .A(\fifo_write/mem[14][4] ), .B(i_wdata[4]), .S0(n1288), .Y(n556) );
  MX2 U1576 ( .A(\fifo_write/mem[14][5] ), .B(i_wdata[5]), .S0(n1288), .Y(n555) );
  MX2 U1577 ( .A(\fifo_write/mem[14][6] ), .B(i_wdata[6]), .S0(n1288), .Y(n554) );
  MX2 U1578 ( .A(\fifo_write/mem[14][7] ), .B(i_wdata[7]), .S0(n1288), .Y(n553) );
  NOR2B U1579 ( .AN(n1373), .B(n1397), .Y(n1398) );
  MX2 U1580 ( .A(\fifo_write/mem[13][0] ), .B(i_wdata[0]), .S0(n1274), .Y(n552) );
  MX2 U1581 ( .A(\fifo_write/mem[13][1] ), .B(i_wdata[1]), .S0(n1274), .Y(n551) );
  MX2 U1582 ( .A(\fifo_write/mem[13][2] ), .B(i_wdata[2]), .S0(n1274), .Y(n550) );
  MX2 U1583 ( .A(\fifo_write/mem[13][3] ), .B(i_wdata[3]), .S0(n1274), .Y(n549) );
  MX2 U1584 ( .A(\fifo_write/mem[13][4] ), .B(i_wdata[4]), .S0(n1274), .Y(n548) );
  MX2 U1585 ( .A(\fifo_write/mem[13][5] ), .B(i_wdata[5]), .S0(n1274), .Y(n547) );
  MX2 U1586 ( .A(\fifo_write/mem[13][6] ), .B(i_wdata[6]), .S0(n1274), .Y(n546) );
  MX2 U1587 ( .A(\fifo_write/mem[13][7] ), .B(i_wdata[7]), .S0(n1274), .Y(n545) );
  NOR2B U1588 ( .AN(n1375), .B(n1397), .Y(n1399) );
  MX2 U1589 ( .A(\fifo_write/mem[12][0] ), .B(i_wdata[0]), .S0(n1276), .Y(n544) );
  MX2 U1590 ( .A(\fifo_write/mem[12][1] ), .B(i_wdata[1]), .S0(n1276), .Y(n543) );
  MX2 U1591 ( .A(\fifo_write/mem[12][2] ), .B(i_wdata[2]), .S0(n1276), .Y(n542) );
  MX2 U1592 ( .A(\fifo_write/mem[12][3] ), .B(i_wdata[3]), .S0(n1276), .Y(n541) );
  MX2 U1593 ( .A(\fifo_write/mem[12][4] ), .B(i_wdata[4]), .S0(n1276), .Y(n540) );
  MX2 U1594 ( .A(\fifo_write/mem[12][5] ), .B(i_wdata[5]), .S0(n1276), .Y(n539) );
  MX2 U1595 ( .A(\fifo_write/mem[12][6] ), .B(i_wdata[6]), .S0(n1276), .Y(n538) );
  MX2 U1596 ( .A(\fifo_write/mem[12][7] ), .B(i_wdata[7]), .S0(n1276), .Y(n537) );
  NOR2B U1597 ( .AN(n1377), .B(n1397), .Y(n1400) );
  MX2 U1598 ( .A(\fifo_write/mem[11][0] ), .B(i_wdata[0]), .S0(n1278), .Y(n536) );
  MX2 U1599 ( .A(\fifo_write/mem[11][1] ), .B(i_wdata[1]), .S0(n1278), .Y(n535) );
  MX2 U1600 ( .A(\fifo_write/mem[11][2] ), .B(i_wdata[2]), .S0(n1278), .Y(n534) );
  MX2 U1601 ( .A(\fifo_write/mem[11][3] ), .B(i_wdata[3]), .S0(n1278), .Y(n533) );
  MX2 U1602 ( .A(\fifo_write/mem[11][4] ), .B(i_wdata[4]), .S0(n1278), .Y(n532) );
  MX2 U1603 ( .A(\fifo_write/mem[11][5] ), .B(i_wdata[5]), .S0(n1278), .Y(n531) );
  MX2 U1604 ( .A(\fifo_write/mem[11][6] ), .B(i_wdata[6]), .S0(n1278), .Y(n530) );
  MX2 U1605 ( .A(\fifo_write/mem[11][7] ), .B(i_wdata[7]), .S0(n1278), .Y(n529) );
  NOR2B U1606 ( .AN(n1379), .B(n1397), .Y(n1401) );
  MX2 U1607 ( .A(\fifo_write/mem[10][0] ), .B(i_wdata[0]), .S0(n1280), .Y(n528) );
  MX2 U1608 ( .A(\fifo_write/mem[10][1] ), .B(i_wdata[1]), .S0(n1280), .Y(n527) );
  MX2 U1609 ( .A(\fifo_write/mem[10][2] ), .B(i_wdata[2]), .S0(n1280), .Y(n526) );
  MX2 U1610 ( .A(\fifo_write/mem[10][3] ), .B(i_wdata[3]), .S0(n1280), .Y(n525) );
  MX2 U1611 ( .A(\fifo_write/mem[10][4] ), .B(i_wdata[4]), .S0(n1280), .Y(n524) );
  MX2 U1612 ( .A(\fifo_write/mem[10][5] ), .B(i_wdata[5]), .S0(n1280), .Y(n523) );
  MX2 U1613 ( .A(\fifo_write/mem[10][6] ), .B(i_wdata[6]), .S0(n1280), .Y(n522) );
  MX2 U1614 ( .A(\fifo_write/mem[10][7] ), .B(i_wdata[7]), .S0(n1280), .Y(n521) );
  NOR2B U1615 ( .AN(n1381), .B(n1397), .Y(n1402) );
  MX2 U1616 ( .A(\fifo_write/mem[9][0] ), .B(i_wdata[0]), .S0(n1266), .Y(n520)
         );
  MX2 U1617 ( .A(\fifo_write/mem[9][1] ), .B(i_wdata[1]), .S0(n1266), .Y(n519)
         );
  MX2 U1618 ( .A(\fifo_write/mem[9][2] ), .B(i_wdata[2]), .S0(n1266), .Y(n518)
         );
  MX2 U1619 ( .A(\fifo_write/mem[9][3] ), .B(i_wdata[3]), .S0(n1266), .Y(n517)
         );
  MX2 U1620 ( .A(\fifo_write/mem[9][4] ), .B(i_wdata[4]), .S0(n1266), .Y(n516)
         );
  MX2 U1621 ( .A(\fifo_write/mem[9][5] ), .B(i_wdata[5]), .S0(n1266), .Y(n515)
         );
  MX2 U1622 ( .A(\fifo_write/mem[9][6] ), .B(i_wdata[6]), .S0(n1266), .Y(n514)
         );
  MX2 U1623 ( .A(\fifo_write/mem[9][7] ), .B(i_wdata[7]), .S0(n1266), .Y(n513)
         );
  NOR2B U1624 ( .AN(n1383), .B(n1397), .Y(n1403) );
  MX2 U1625 ( .A(\fifo_write/mem[8][0] ), .B(i_wdata[0]), .S0(n1268), .Y(n512)
         );
  MX2 U1626 ( .A(\fifo_write/mem[8][1] ), .B(i_wdata[1]), .S0(n1268), .Y(n511)
         );
  MX2 U1627 ( .A(\fifo_write/mem[8][2] ), .B(i_wdata[2]), .S0(n1268), .Y(n510)
         );
  MX2 U1628 ( .A(\fifo_write/mem[8][3] ), .B(i_wdata[3]), .S0(n1268), .Y(n509)
         );
  MX2 U1629 ( .A(\fifo_write/mem[8][4] ), .B(i_wdata[4]), .S0(n1268), .Y(n508)
         );
  MX2 U1630 ( .A(\fifo_write/mem[8][5] ), .B(i_wdata[5]), .S0(n1268), .Y(n507)
         );
  MX2 U1631 ( .A(\fifo_write/mem[8][6] ), .B(i_wdata[6]), .S0(n1268), .Y(n506)
         );
  MX2 U1632 ( .A(\fifo_write/mem[8][7] ), .B(i_wdata[7]), .S0(n1268), .Y(n505)
         );
  NOR2B U1633 ( .AN(n1385), .B(n1397), .Y(n1404) );
  NAND3B U1634 ( .AN(\fifo_write/waddr[4] ), .B(n1386), .C(
        \fifo_write/waddr[3] ), .Y(n1397) );
  MX2 U1635 ( .A(\fifo_write/mem[7][0] ), .B(i_wdata[0]), .S0(n1270), .Y(n504)
         );
  MX2 U1636 ( .A(\fifo_write/mem[7][1] ), .B(i_wdata[1]), .S0(n1270), .Y(n503)
         );
  MX2 U1637 ( .A(\fifo_write/mem[7][2] ), .B(i_wdata[2]), .S0(n1270), .Y(n502)
         );
  MX2 U1638 ( .A(\fifo_write/mem[7][3] ), .B(i_wdata[3]), .S0(n1270), .Y(n501)
         );
  MX2 U1639 ( .A(\fifo_write/mem[7][4] ), .B(i_wdata[4]), .S0(n1270), .Y(n500)
         );
  MX2 U1640 ( .A(\fifo_write/mem[7][5] ), .B(i_wdata[5]), .S0(n1270), .Y(n499)
         );
  MX2 U1641 ( .A(\fifo_write/mem[7][6] ), .B(i_wdata[6]), .S0(n1270), .Y(n498)
         );
  MX2 U1642 ( .A(\fifo_write/mem[7][7] ), .B(i_wdata[7]), .S0(n1270), .Y(n497)
         );
  NOR2B U1643 ( .AN(n1370), .B(n1406), .Y(n1405) );
  NOR3B U1644 ( .AN(\fifo_write/waddr[2] ), .B(n1407), .C(n1408), .Y(n1370) );
  MX2 U1645 ( .A(\fifo_write/mem[6][0] ), .B(i_wdata[0]), .S0(n1272), .Y(n496)
         );
  MX2 U1646 ( .A(\fifo_write/mem[6][1] ), .B(i_wdata[1]), .S0(n1272), .Y(n495)
         );
  MX2 U1647 ( .A(\fifo_write/mem[6][2] ), .B(i_wdata[2]), .S0(n1272), .Y(n494)
         );
  MX2 U1648 ( .A(\fifo_write/mem[6][3] ), .B(i_wdata[3]), .S0(n1272), .Y(n493)
         );
  MX2 U1649 ( .A(\fifo_write/mem[6][4] ), .B(i_wdata[4]), .S0(n1272), .Y(n492)
         );
  MX2 U1650 ( .A(\fifo_write/mem[6][5] ), .B(i_wdata[5]), .S0(n1272), .Y(n491)
         );
  MX2 U1651 ( .A(\fifo_write/mem[6][6] ), .B(i_wdata[6]), .S0(n1272), .Y(n490)
         );
  MX2 U1652 ( .A(\fifo_write/mem[6][7] ), .B(i_wdata[7]), .S0(n1272), .Y(n489)
         );
  NOR2B U1653 ( .AN(n1373), .B(n1406), .Y(n1409) );
  NOR3B U1654 ( .AN(\fifo_write/waddr[2] ), .B(\fifo_write/waddr[0] ), .C(
        n1408), .Y(n1373) );
  MX2 U1655 ( .A(\fifo_write/mem[5][0] ), .B(i_wdata[0]), .S0(n1262), .Y(n488)
         );
  MX2 U1656 ( .A(\fifo_write/mem[5][1] ), .B(i_wdata[1]), .S0(n1262), .Y(n487)
         );
  MX2 U1657 ( .A(\fifo_write/mem[5][2] ), .B(i_wdata[2]), .S0(n1262), .Y(n486)
         );
  MX2 U1658 ( .A(\fifo_write/mem[5][3] ), .B(i_wdata[3]), .S0(n1262), .Y(n485)
         );
  MX2 U1659 ( .A(\fifo_write/mem[5][4] ), .B(i_wdata[4]), .S0(n1262), .Y(n484)
         );
  MX2 U1660 ( .A(\fifo_write/mem[5][5] ), .B(i_wdata[5]), .S0(n1262), .Y(n483)
         );
  MX2 U1661 ( .A(\fifo_write/mem[5][6] ), .B(i_wdata[6]), .S0(n1262), .Y(n482)
         );
  MX2 U1662 ( .A(\fifo_write/mem[5][7] ), .B(i_wdata[7]), .S0(n1262), .Y(n481)
         );
  NOR2B U1663 ( .AN(n1375), .B(n1406), .Y(n1410) );
  NOR3B U1664 ( .AN(\fifo_write/waddr[2] ), .B(\fifo_write/waddr[1] ), .C(
        n1407), .Y(n1375) );
  MX2 U1665 ( .A(\fifo_write/mem[4][0] ), .B(i_wdata[0]), .S0(n1264), .Y(n480)
         );
  MX2 U1666 ( .A(\fifo_write/mem[4][1] ), .B(i_wdata[1]), .S0(n1264), .Y(n479)
         );
  MX2 U1667 ( .A(\fifo_write/mem[4][2] ), .B(i_wdata[2]), .S0(n1264), .Y(n478)
         );
  MX2 U1668 ( .A(\fifo_write/mem[4][3] ), .B(i_wdata[3]), .S0(n1264), .Y(n477)
         );
  MX2 U1669 ( .A(\fifo_write/mem[4][4] ), .B(i_wdata[4]), .S0(n1264), .Y(n476)
         );
  MX2 U1670 ( .A(\fifo_write/mem[4][5] ), .B(i_wdata[5]), .S0(n1264), .Y(n475)
         );
  MX2 U1671 ( .A(\fifo_write/mem[4][6] ), .B(i_wdata[6]), .S0(n1264), .Y(n474)
         );
  MX2 U1672 ( .A(\fifo_write/mem[4][7] ), .B(i_wdata[7]), .S0(n1264), .Y(n473)
         );
  NOR2B U1673 ( .AN(n1377), .B(n1406), .Y(n1411) );
  NOR3B U1674 ( .AN(\fifo_write/waddr[2] ), .B(\fifo_write/waddr[0] ), .C(
        \fifo_write/waddr[1] ), .Y(n1377) );
  MX2 U1675 ( .A(\fifo_write/mem[3][0] ), .B(i_wdata[0]), .S0(n1258), .Y(n472)
         );
  MX2 U1676 ( .A(\fifo_write/mem[3][1] ), .B(i_wdata[1]), .S0(n1258), .Y(n471)
         );
  MX2 U1677 ( .A(\fifo_write/mem[3][2] ), .B(i_wdata[2]), .S0(n1258), .Y(n470)
         );
  MX2 U1678 ( .A(\fifo_write/mem[3][3] ), .B(i_wdata[3]), .S0(n1258), .Y(n469)
         );
  MX2 U1679 ( .A(\fifo_write/mem[3][4] ), .B(i_wdata[4]), .S0(n1258), .Y(n468)
         );
  MX2 U1680 ( .A(\fifo_write/mem[3][5] ), .B(i_wdata[5]), .S0(n1258), .Y(n467)
         );
  MX2 U1681 ( .A(\fifo_write/mem[3][6] ), .B(i_wdata[6]), .S0(n1258), .Y(n466)
         );
  MX2 U1682 ( .A(\fifo_write/mem[3][7] ), .B(i_wdata[7]), .S0(n1258), .Y(n465)
         );
  NOR2B U1683 ( .AN(n1379), .B(n1406), .Y(n1412) );
  NOR3 U1684 ( .A(\fifo_write/waddr[2] ), .B(n1407), .C(n1408), .Y(n1379) );
  MX2 U1685 ( .A(\fifo_write/mem[2][0] ), .B(i_wdata[0]), .S0(n1260), .Y(n464)
         );
  MX2 U1686 ( .A(\fifo_write/mem[2][1] ), .B(i_wdata[1]), .S0(n1260), .Y(n463)
         );
  MX2 U1687 ( .A(\fifo_write/mem[2][2] ), .B(i_wdata[2]), .S0(n1260), .Y(n462)
         );
  MX2 U1688 ( .A(\fifo_write/mem[2][3] ), .B(i_wdata[3]), .S0(n1260), .Y(n461)
         );
  MX2 U1689 ( .A(\fifo_write/mem[2][4] ), .B(i_wdata[4]), .S0(n1260), .Y(n460)
         );
  MX2 U1690 ( .A(\fifo_write/mem[2][5] ), .B(i_wdata[5]), .S0(n1260), .Y(n459)
         );
  MX2 U1691 ( .A(\fifo_write/mem[2][6] ), .B(i_wdata[6]), .S0(n1260), .Y(n458)
         );
  MX2 U1692 ( .A(\fifo_write/mem[2][7] ), .B(i_wdata[7]), .S0(n1260), .Y(n457)
         );
  NOR2B U1693 ( .AN(n1381), .B(n1406), .Y(n1413) );
  NOR3 U1694 ( .A(\fifo_write/waddr[2] ), .B(\fifo_write/waddr[0] ), .C(n1408), 
        .Y(n1381) );
  MX2 U1695 ( .A(\fifo_write/mem[1][0] ), .B(i_wdata[0]), .S0(n1254), .Y(n456)
         );
  MX2 U1696 ( .A(\fifo_write/mem[1][1] ), .B(i_wdata[1]), .S0(n1254), .Y(n455)
         );
  MX2 U1697 ( .A(\fifo_write/mem[1][2] ), .B(i_wdata[2]), .S0(n1254), .Y(n454)
         );
  MX2 U1698 ( .A(\fifo_write/mem[1][3] ), .B(i_wdata[3]), .S0(n1254), .Y(n453)
         );
  MX2 U1699 ( .A(\fifo_write/mem[1][4] ), .B(i_wdata[4]), .S0(n1254), .Y(n452)
         );
  MX2 U1700 ( .A(\fifo_write/mem[1][5] ), .B(i_wdata[5]), .S0(n1254), .Y(n451)
         );
  MX2 U1701 ( .A(\fifo_write/mem[1][6] ), .B(i_wdata[6]), .S0(n1254), .Y(n450)
         );
  MX2 U1702 ( .A(\fifo_write/mem[1][7] ), .B(i_wdata[7]), .S0(n1254), .Y(n449)
         );
  NOR2B U1703 ( .AN(n1383), .B(n1406), .Y(n1414) );
  NOR2B U1704 ( .AN(n1415), .B(n1407), .Y(n1383) );
  MX2 U1705 ( .A(\fifo_write/mem[0][0] ), .B(i_wdata[0]), .S0(n1256), .Y(n448)
         );
  MX2 U1706 ( .A(\fifo_write/mem[0][1] ), .B(i_wdata[1]), .S0(n1256), .Y(n447)
         );
  MX2 U1707 ( .A(\fifo_write/mem[0][2] ), .B(i_wdata[2]), .S0(n1256), .Y(n446)
         );
  MX2 U1708 ( .A(\fifo_write/mem[0][3] ), .B(i_wdata[3]), .S0(n1256), .Y(n445)
         );
  MX2 U1709 ( .A(\fifo_write/mem[0][4] ), .B(i_wdata[4]), .S0(n1256), .Y(n444)
         );
  MX2 U1710 ( .A(\fifo_write/mem[0][5] ), .B(i_wdata[5]), .S0(n1256), .Y(n443)
         );
  MX2 U1711 ( .A(\fifo_write/mem[0][6] ), .B(i_wdata[6]), .S0(n1256), .Y(n442)
         );
  MX2 U1712 ( .A(\fifo_write/mem[0][7] ), .B(i_wdata[7]), .S0(n1256), .Y(n441)
         );
  NOR2B U1713 ( .AN(n1385), .B(n1406), .Y(n1416) );
  INV U1714 ( .A(n1417), .Y(n1406) );
  NOR3B U1715 ( .AN(n1386), .B(\fifo_write/waddr[4] ), .C(
        \fifo_write/waddr[3] ), .Y(n1417) );
  NOR2B U1716 ( .AN(n1415), .B(\fifo_write/waddr[0] ), .Y(n1385) );
  NOR2 U1717 ( .A(\fifo_write/waddr[2] ), .B(\fifo_write/waddr[1] ), .Y(n1415)
         );
  MX2 U1718 ( .A(\fifo_read/mem[31][0] ), .B(wdata_to_fifo[0]), .S0(n1250), 
        .Y(n440) );
  MX2 U1719 ( .A(\fifo_read/mem[31][1] ), .B(wdata_to_fifo[1]), .S0(n1250), 
        .Y(n439) );
  MX2 U1720 ( .A(\fifo_read/mem[31][2] ), .B(n1328), .S0(n1250), .Y(n438) );
  MX2 U1721 ( .A(\fifo_read/mem[31][3] ), .B(n1326), .S0(n1250), .Y(n437) );
  MX2 U1722 ( .A(\fifo_read/mem[31][4] ), .B(n1324), .S0(n1250), .Y(n436) );
  MX2 U1723 ( .A(\fifo_read/mem[31][5] ), .B(n1322), .S0(n1250), .Y(n435) );
  MX2 U1724 ( .A(\fifo_read/mem[31][6] ), .B(n1336), .S0(n1250), .Y(n434) );
  MX2 U1725 ( .A(\fifo_read/mem[31][7] ), .B(wdata_to_fifo[7]), .S0(n1250), 
        .Y(n433) );
  NOR2B U1726 ( .AN(n1419), .B(n1420), .Y(n1418) );
  MX2 U1727 ( .A(\fifo_read/mem[30][0] ), .B(n1316), .S0(n1252), .Y(n432) );
  MX2 U1728 ( .A(\fifo_read/mem[30][1] ), .B(n1314), .S0(n1252), .Y(n431) );
  MX2 U1729 ( .A(\fifo_read/mem[30][2] ), .B(n1328), .S0(n1252), .Y(n430) );
  MX2 U1730 ( .A(\fifo_read/mem[30][3] ), .B(n1326), .S0(n1252), .Y(n429) );
  MX2 U1731 ( .A(\fifo_read/mem[30][4] ), .B(n1324), .S0(n1252), .Y(n428) );
  MX2 U1732 ( .A(\fifo_read/mem[30][5] ), .B(n1322), .S0(n1252), .Y(n427) );
  MX2 U1733 ( .A(\fifo_read/mem[30][6] ), .B(n1336), .S0(n1252), .Y(n426) );
  MX2 U1734 ( .A(\fifo_read/mem[30][7] ), .B(n1334), .S0(n1252), .Y(n425) );
  NOR2B U1735 ( .AN(n1422), .B(n1420), .Y(n1421) );
  MX2 U1736 ( .A(\fifo_read/mem[29][0] ), .B(wdata_to_fifo[0]), .S0(n1246), 
        .Y(n424) );
  MX2 U1737 ( .A(\fifo_read/mem[29][1] ), .B(wdata_to_fifo[1]), .S0(n1246), 
        .Y(n423) );
  MX2 U1738 ( .A(\fifo_read/mem[29][2] ), .B(wdata_to_fifo[2]), .S0(n1246), 
        .Y(n422) );
  MX2 U1739 ( .A(\fifo_read/mem[29][3] ), .B(wdata_to_fifo[3]), .S0(n1246), 
        .Y(n421) );
  MX2 U1740 ( .A(\fifo_read/mem[29][4] ), .B(wdata_to_fifo[4]), .S0(n1246), 
        .Y(n420) );
  MX2 U1741 ( .A(\fifo_read/mem[29][5] ), .B(wdata_to_fifo[5]), .S0(n1246), 
        .Y(n419) );
  MX2 U1742 ( .A(\fifo_read/mem[29][6] ), .B(wdata_to_fifo[6]), .S0(n1246), 
        .Y(n418) );
  MX2 U1743 ( .A(\fifo_read/mem[29][7] ), .B(wdata_to_fifo[7]), .S0(n1246), 
        .Y(n417) );
  NOR2B U1744 ( .AN(n1424), .B(n1420), .Y(n1423) );
  MX2 U1745 ( .A(\fifo_read/mem[28][0] ), .B(n1316), .S0(n1248), .Y(n416) );
  MX2 U1746 ( .A(\fifo_read/mem[28][1] ), .B(n1314), .S0(n1248), .Y(n415) );
  MX2 U1747 ( .A(\fifo_read/mem[28][2] ), .B(n1328), .S0(n1248), .Y(n414) );
  MX2 U1748 ( .A(\fifo_read/mem[28][3] ), .B(n1326), .S0(n1248), .Y(n413) );
  MX2 U1749 ( .A(\fifo_read/mem[28][4] ), .B(n1324), .S0(n1248), .Y(n412) );
  MX2 U1750 ( .A(\fifo_read/mem[28][5] ), .B(n1322), .S0(n1248), .Y(n411) );
  MX2 U1751 ( .A(\fifo_read/mem[28][6] ), .B(n1336), .S0(n1248), .Y(n410) );
  MX2 U1752 ( .A(\fifo_read/mem[28][7] ), .B(n1334), .S0(n1248), .Y(n409) );
  NOR2B U1753 ( .AN(n1426), .B(n1420), .Y(n1425) );
  MX2 U1754 ( .A(\fifo_read/mem[27][0] ), .B(wdata_to_fifo[0]), .S0(n1242), 
        .Y(n408) );
  MX2 U1755 ( .A(\fifo_read/mem[27][1] ), .B(wdata_to_fifo[1]), .S0(n1242), 
        .Y(n407) );
  MX2 U1756 ( .A(\fifo_read/mem[27][2] ), .B(wdata_to_fifo[2]), .S0(n1242), 
        .Y(n406) );
  MX2 U1757 ( .A(\fifo_read/mem[27][3] ), .B(wdata_to_fifo[3]), .S0(n1242), 
        .Y(n405) );
  MX2 U1758 ( .A(\fifo_read/mem[27][4] ), .B(wdata_to_fifo[4]), .S0(n1242), 
        .Y(n404) );
  MX2 U1759 ( .A(\fifo_read/mem[27][5] ), .B(wdata_to_fifo[5]), .S0(n1242), 
        .Y(n403) );
  MX2 U1760 ( .A(\fifo_read/mem[27][6] ), .B(wdata_to_fifo[6]), .S0(n1242), 
        .Y(n402) );
  MX2 U1761 ( .A(\fifo_read/mem[27][7] ), .B(wdata_to_fifo[7]), .S0(n1242), 
        .Y(n401) );
  NOR2B U1762 ( .AN(n1428), .B(n1420), .Y(n1427) );
  MX2 U1763 ( .A(\fifo_read/mem[26][0] ), .B(n1316), .S0(n1244), .Y(n400) );
  MX2 U1764 ( .A(\fifo_read/mem[26][1] ), .B(n1314), .S0(n1244), .Y(n399) );
  MX2 U1765 ( .A(\fifo_read/mem[26][2] ), .B(n1328), .S0(n1244), .Y(n398) );
  MX2 U1766 ( .A(\fifo_read/mem[26][3] ), .B(n1326), .S0(n1244), .Y(n397) );
  MX2 U1767 ( .A(\fifo_read/mem[26][4] ), .B(n1324), .S0(n1244), .Y(n396) );
  MX2 U1768 ( .A(\fifo_read/mem[26][5] ), .B(n1322), .S0(n1244), .Y(n395) );
  MX2 U1769 ( .A(\fifo_read/mem[26][6] ), .B(n1336), .S0(n1244), .Y(n394) );
  MX2 U1770 ( .A(\fifo_read/mem[26][7] ), .B(n1334), .S0(n1244), .Y(n393) );
  NOR2B U1771 ( .AN(n1430), .B(n1420), .Y(n1429) );
  MX2 U1772 ( .A(\fifo_read/mem[25][0] ), .B(wdata_to_fifo[0]), .S0(n1238), 
        .Y(n392) );
  MX2 U1773 ( .A(\fifo_read/mem[25][1] ), .B(wdata_to_fifo[1]), .S0(n1238), 
        .Y(n391) );
  MX2 U1774 ( .A(\fifo_read/mem[25][2] ), .B(wdata_to_fifo[2]), .S0(n1238), 
        .Y(n390) );
  MX2 U1775 ( .A(\fifo_read/mem[25][3] ), .B(wdata_to_fifo[3]), .S0(n1238), 
        .Y(n389) );
  MX2 U1776 ( .A(\fifo_read/mem[25][4] ), .B(wdata_to_fifo[4]), .S0(n1238), 
        .Y(n388) );
  MX2 U1777 ( .A(\fifo_read/mem[25][5] ), .B(wdata_to_fifo[5]), .S0(n1238), 
        .Y(n387) );
  MX2 U1778 ( .A(\fifo_read/mem[25][6] ), .B(wdata_to_fifo[6]), .S0(n1238), 
        .Y(n386) );
  MX2 U1779 ( .A(\fifo_read/mem[25][7] ), .B(wdata_to_fifo[7]), .S0(n1238), 
        .Y(n385) );
  NOR2B U1780 ( .AN(n1432), .B(n1420), .Y(n1431) );
  MX2 U1781 ( .A(\fifo_read/mem[24][0] ), .B(n1316), .S0(n1240), .Y(n384) );
  MX2 U1782 ( .A(\fifo_read/mem[24][1] ), .B(n1314), .S0(n1240), .Y(n383) );
  MX2 U1783 ( .A(\fifo_read/mem[24][2] ), .B(n1328), .S0(n1240), .Y(n382) );
  MX2 U1784 ( .A(\fifo_read/mem[24][3] ), .B(n1326), .S0(n1240), .Y(n381) );
  MX2 U1785 ( .A(\fifo_read/mem[24][4] ), .B(n1324), .S0(n1240), .Y(n380) );
  MX2 U1786 ( .A(\fifo_read/mem[24][5] ), .B(n1322), .S0(n1240), .Y(n379) );
  MX2 U1787 ( .A(\fifo_read/mem[24][6] ), .B(n1336), .S0(n1240), .Y(n378) );
  MX2 U1788 ( .A(\fifo_read/mem[24][7] ), .B(n1334), .S0(n1240), .Y(n377) );
  NOR2B U1789 ( .AN(n1434), .B(n1420), .Y(n1433) );
  NAND3 U1790 ( .A(n1435), .B(\fifo_read/waddr[4] ), .C(\fifo_read/waddr[3] ), 
        .Y(n1420) );
  MX2 U1791 ( .A(\fifo_read/mem[23][0] ), .B(wdata_to_fifo[0]), .S0(n1234), 
        .Y(n376) );
  MX2 U1792 ( .A(\fifo_read/mem[23][1] ), .B(wdata_to_fifo[1]), .S0(n1234), 
        .Y(n375) );
  MX2 U1793 ( .A(\fifo_read/mem[23][2] ), .B(wdata_to_fifo[2]), .S0(n1234), 
        .Y(n374) );
  MX2 U1794 ( .A(\fifo_read/mem[23][3] ), .B(wdata_to_fifo[3]), .S0(n1234), 
        .Y(n373) );
  MX2 U1795 ( .A(\fifo_read/mem[23][4] ), .B(wdata_to_fifo[4]), .S0(n1234), 
        .Y(n372) );
  MX2 U1796 ( .A(\fifo_read/mem[23][5] ), .B(wdata_to_fifo[5]), .S0(n1234), 
        .Y(n371) );
  MX2 U1797 ( .A(\fifo_read/mem[23][6] ), .B(wdata_to_fifo[6]), .S0(n1234), 
        .Y(n370) );
  MX2 U1798 ( .A(\fifo_read/mem[23][7] ), .B(wdata_to_fifo[7]), .S0(n1234), 
        .Y(n369) );
  NOR2B U1799 ( .AN(n1419), .B(n1437), .Y(n1436) );
  MX2 U1800 ( .A(\fifo_read/mem[22][0] ), .B(n1316), .S0(n1236), .Y(n368) );
  MX2 U1801 ( .A(\fifo_read/mem[22][1] ), .B(n1314), .S0(n1236), .Y(n367) );
  MX2 U1802 ( .A(\fifo_read/mem[22][2] ), .B(n1328), .S0(n1236), .Y(n366) );
  MX2 U1803 ( .A(\fifo_read/mem[22][3] ), .B(n1326), .S0(n1236), .Y(n365) );
  MX2 U1804 ( .A(\fifo_read/mem[22][4] ), .B(n1324), .S0(n1236), .Y(n364) );
  MX2 U1805 ( .A(\fifo_read/mem[22][5] ), .B(n1322), .S0(n1236), .Y(n363) );
  MX2 U1806 ( .A(\fifo_read/mem[22][6] ), .B(n1336), .S0(n1236), .Y(n362) );
  MX2 U1807 ( .A(\fifo_read/mem[22][7] ), .B(n1334), .S0(n1236), .Y(n361) );
  NOR2B U1808 ( .AN(n1422), .B(n1437), .Y(n1438) );
  MX2 U1809 ( .A(\fifo_read/mem[21][0] ), .B(wdata_to_fifo[0]), .S0(n1230), 
        .Y(n360) );
  MX2 U1810 ( .A(\fifo_read/mem[21][1] ), .B(wdata_to_fifo[1]), .S0(n1230), 
        .Y(n359) );
  MX2 U1811 ( .A(\fifo_read/mem[21][2] ), .B(wdata_to_fifo[2]), .S0(n1230), 
        .Y(n358) );
  MX2 U1812 ( .A(\fifo_read/mem[21][3] ), .B(wdata_to_fifo[3]), .S0(n1230), 
        .Y(n357) );
  MX2 U1813 ( .A(\fifo_read/mem[21][4] ), .B(wdata_to_fifo[4]), .S0(n1230), 
        .Y(n356) );
  MX2 U1814 ( .A(\fifo_read/mem[21][5] ), .B(wdata_to_fifo[5]), .S0(n1230), 
        .Y(n355) );
  MX2 U1815 ( .A(\fifo_read/mem[21][6] ), .B(wdata_to_fifo[6]), .S0(n1230), 
        .Y(n354) );
  MX2 U1816 ( .A(\fifo_read/mem[21][7] ), .B(wdata_to_fifo[7]), .S0(n1230), 
        .Y(n353) );
  NOR2B U1817 ( .AN(n1424), .B(n1437), .Y(n1439) );
  MX2 U1818 ( .A(\fifo_read/mem[20][0] ), .B(n1316), .S0(n1232), .Y(n352) );
  MX2 U1819 ( .A(\fifo_read/mem[20][1] ), .B(n1314), .S0(n1232), .Y(n351) );
  MX2 U1820 ( .A(\fifo_read/mem[20][2] ), .B(n1328), .S0(n1232), .Y(n350) );
  MX2 U1821 ( .A(\fifo_read/mem[20][3] ), .B(n1326), .S0(n1232), .Y(n349) );
  MX2 U1822 ( .A(\fifo_read/mem[20][4] ), .B(n1324), .S0(n1232), .Y(n348) );
  MX2 U1823 ( .A(\fifo_read/mem[20][5] ), .B(n1322), .S0(n1232), .Y(n347) );
  MX2 U1824 ( .A(\fifo_read/mem[20][6] ), .B(n1336), .S0(n1232), .Y(n346) );
  MX2 U1825 ( .A(\fifo_read/mem[20][7] ), .B(n1334), .S0(n1232), .Y(n345) );
  NOR2B U1826 ( .AN(n1426), .B(n1437), .Y(n1440) );
  MX2 U1827 ( .A(\fifo_read/mem[19][0] ), .B(wdata_to_fifo[0]), .S0(n1226), 
        .Y(n344) );
  MX2 U1828 ( .A(\fifo_read/mem[19][1] ), .B(wdata_to_fifo[1]), .S0(n1226), 
        .Y(n343) );
  MX2 U1829 ( .A(\fifo_read/mem[19][2] ), .B(wdata_to_fifo[2]), .S0(n1226), 
        .Y(n342) );
  MX2 U1830 ( .A(\fifo_read/mem[19][3] ), .B(wdata_to_fifo[3]), .S0(n1226), 
        .Y(n341) );
  MX2 U1831 ( .A(\fifo_read/mem[19][4] ), .B(wdata_to_fifo[4]), .S0(n1226), 
        .Y(n340) );
  MX2 U1832 ( .A(\fifo_read/mem[19][5] ), .B(wdata_to_fifo[5]), .S0(n1226), 
        .Y(n339) );
  MX2 U1833 ( .A(\fifo_read/mem[19][6] ), .B(wdata_to_fifo[6]), .S0(n1226), 
        .Y(n338) );
  MX2 U1834 ( .A(\fifo_read/mem[19][7] ), .B(wdata_to_fifo[7]), .S0(n1226), 
        .Y(n337) );
  NOR2B U1835 ( .AN(n1428), .B(n1437), .Y(n1441) );
  MX2 U1836 ( .A(\fifo_read/mem[18][0] ), .B(n1316), .S0(n1228), .Y(n336) );
  MX2 U1837 ( .A(\fifo_read/mem[18][1] ), .B(n1314), .S0(n1228), .Y(n335) );
  MX2 U1838 ( .A(\fifo_read/mem[18][2] ), .B(n1328), .S0(n1228), .Y(n334) );
  MX2 U1839 ( .A(\fifo_read/mem[18][3] ), .B(n1326), .S0(n1228), .Y(n333) );
  MX2 U1840 ( .A(\fifo_read/mem[18][4] ), .B(n1324), .S0(n1228), .Y(n332) );
  MX2 U1841 ( .A(\fifo_read/mem[18][5] ), .B(n1322), .S0(n1228), .Y(n331) );
  MX2 U1842 ( .A(\fifo_read/mem[18][6] ), .B(n1336), .S0(n1228), .Y(n330) );
  MX2 U1843 ( .A(\fifo_read/mem[18][7] ), .B(n1334), .S0(n1228), .Y(n329) );
  NOR2B U1844 ( .AN(n1430), .B(n1437), .Y(n1442) );
  MX2 U1845 ( .A(\fifo_read/mem[17][0] ), .B(wdata_to_fifo[0]), .S0(n1222), 
        .Y(n328) );
  MX2 U1846 ( .A(\fifo_read/mem[17][1] ), .B(wdata_to_fifo[1]), .S0(n1222), 
        .Y(n327) );
  MX2 U1847 ( .A(\fifo_read/mem[17][2] ), .B(wdata_to_fifo[2]), .S0(n1222), 
        .Y(n326) );
  MX2 U1848 ( .A(\fifo_read/mem[17][3] ), .B(wdata_to_fifo[3]), .S0(n1222), 
        .Y(n325) );
  MX2 U1849 ( .A(\fifo_read/mem[17][4] ), .B(wdata_to_fifo[4]), .S0(n1222), 
        .Y(n324) );
  MX2 U1850 ( .A(\fifo_read/mem[17][5] ), .B(wdata_to_fifo[5]), .S0(n1222), 
        .Y(n323) );
  MX2 U1851 ( .A(\fifo_read/mem[17][6] ), .B(wdata_to_fifo[6]), .S0(n1222), 
        .Y(n322) );
  MX2 U1852 ( .A(\fifo_read/mem[17][7] ), .B(wdata_to_fifo[7]), .S0(n1222), 
        .Y(n321) );
  NOR2B U1853 ( .AN(n1432), .B(n1437), .Y(n1443) );
  MX2 U1854 ( .A(\fifo_read/mem[16][0] ), .B(n1316), .S0(n1224), .Y(n320) );
  MX2 U1855 ( .A(\fifo_read/mem[16][1] ), .B(n1314), .S0(n1224), .Y(n319) );
  MX2 U1856 ( .A(\fifo_read/mem[16][2] ), .B(n1328), .S0(n1224), .Y(n318) );
  MX2 U1857 ( .A(\fifo_read/mem[16][3] ), .B(n1326), .S0(n1224), .Y(n317) );
  MX2 U1858 ( .A(\fifo_read/mem[16][4] ), .B(n1324), .S0(n1224), .Y(n316) );
  MX2 U1859 ( .A(\fifo_read/mem[16][5] ), .B(n1322), .S0(n1224), .Y(n315) );
  MX2 U1860 ( .A(\fifo_read/mem[16][6] ), .B(n1336), .S0(n1224), .Y(n314) );
  MX2 U1861 ( .A(\fifo_read/mem[16][7] ), .B(n1334), .S0(n1224), .Y(n313) );
  NOR2B U1862 ( .AN(n1434), .B(n1437), .Y(n1444) );
  NAND3B U1863 ( .AN(\fifo_read/waddr[3] ), .B(\fifo_read/waddr[4] ), .C(n1435), .Y(n1437) );
  MX2 U1864 ( .A(\fifo_read/mem[15][0] ), .B(wdata_to_fifo[0]), .S0(n1218), 
        .Y(n312) );
  MX2 U1865 ( .A(\fifo_read/mem[15][1] ), .B(wdata_to_fifo[1]), .S0(n1218), 
        .Y(n311) );
  MX2 U1866 ( .A(\fifo_read/mem[15][2] ), .B(wdata_to_fifo[2]), .S0(n1218), 
        .Y(n310) );
  MX2 U1867 ( .A(\fifo_read/mem[15][3] ), .B(wdata_to_fifo[3]), .S0(n1218), 
        .Y(n309) );
  MX2 U1868 ( .A(\fifo_read/mem[15][4] ), .B(wdata_to_fifo[4]), .S0(n1218), 
        .Y(n308) );
  MX2 U1869 ( .A(\fifo_read/mem[15][5] ), .B(wdata_to_fifo[5]), .S0(n1218), 
        .Y(n307) );
  MX2 U1870 ( .A(\fifo_read/mem[15][6] ), .B(wdata_to_fifo[6]), .S0(n1218), 
        .Y(n306) );
  MX2 U1871 ( .A(\fifo_read/mem[15][7] ), .B(wdata_to_fifo[7]), .S0(n1218), 
        .Y(n305) );
  NOR2B U1872 ( .AN(n1419), .B(n1446), .Y(n1445) );
  MX2 U1873 ( .A(\fifo_read/mem[14][0] ), .B(n1316), .S0(n1220), .Y(n304) );
  MX2 U1874 ( .A(\fifo_read/mem[14][1] ), .B(n1314), .S0(n1220), .Y(n303) );
  MX2 U1875 ( .A(\fifo_read/mem[14][2] ), .B(n1328), .S0(n1220), .Y(n302) );
  MX2 U1876 ( .A(\fifo_read/mem[14][3] ), .B(n1326), .S0(n1220), .Y(n301) );
  MX2 U1877 ( .A(\fifo_read/mem[14][4] ), .B(n1324), .S0(n1220), .Y(n300) );
  MX2 U1878 ( .A(\fifo_read/mem[14][5] ), .B(n1322), .S0(n1220), .Y(n299) );
  MX2 U1879 ( .A(\fifo_read/mem[14][6] ), .B(n1336), .S0(n1220), .Y(n298) );
  MX2 U1880 ( .A(\fifo_read/mem[14][7] ), .B(n1334), .S0(n1220), .Y(n297) );
  NOR2B U1881 ( .AN(n1422), .B(n1446), .Y(n1447) );
  MX2 U1882 ( .A(\fifo_read/mem[13][0] ), .B(wdata_to_fifo[0]), .S0(n1214), 
        .Y(n296) );
  MX2 U1883 ( .A(\fifo_read/mem[13][1] ), .B(wdata_to_fifo[1]), .S0(n1214), 
        .Y(n295) );
  MX2 U1884 ( .A(\fifo_read/mem[13][2] ), .B(wdata_to_fifo[2]), .S0(n1214), 
        .Y(n294) );
  MX2 U1885 ( .A(\fifo_read/mem[13][3] ), .B(wdata_to_fifo[3]), .S0(n1214), 
        .Y(n293) );
  MX2 U1886 ( .A(\fifo_read/mem[13][4] ), .B(wdata_to_fifo[4]), .S0(n1214), 
        .Y(n292) );
  MX2 U1887 ( .A(\fifo_read/mem[13][5] ), .B(wdata_to_fifo[5]), .S0(n1214), 
        .Y(n291) );
  MX2 U1888 ( .A(\fifo_read/mem[13][6] ), .B(wdata_to_fifo[6]), .S0(n1214), 
        .Y(n290) );
  MX2 U1889 ( .A(\fifo_read/mem[13][7] ), .B(wdata_to_fifo[7]), .S0(n1214), 
        .Y(n289) );
  NOR2B U1890 ( .AN(n1424), .B(n1446), .Y(n1448) );
  MX2 U1891 ( .A(\fifo_read/mem[12][0] ), .B(n1316), .S0(n1216), .Y(n288) );
  MX2 U1892 ( .A(\fifo_read/mem[12][1] ), .B(n1314), .S0(n1216), .Y(n287) );
  MX2 U1893 ( .A(\fifo_read/mem[12][2] ), .B(n1328), .S0(n1216), .Y(n286) );
  MX2 U1894 ( .A(\fifo_read/mem[12][3] ), .B(n1326), .S0(n1216), .Y(n285) );
  MX2 U1895 ( .A(\fifo_read/mem[12][4] ), .B(n1324), .S0(n1216), .Y(n284) );
  MX2 U1896 ( .A(\fifo_read/mem[12][5] ), .B(n1322), .S0(n1216), .Y(n283) );
  MX2 U1897 ( .A(\fifo_read/mem[12][6] ), .B(n1336), .S0(n1216), .Y(n282) );
  MX2 U1898 ( .A(\fifo_read/mem[12][7] ), .B(n1334), .S0(n1216), .Y(n281) );
  NOR2B U1899 ( .AN(n1426), .B(n1446), .Y(n1449) );
  MX2 U1900 ( .A(\fifo_read/mem[11][0] ), .B(wdata_to_fifo[0]), .S0(n1210), 
        .Y(n280) );
  MX2 U1901 ( .A(\fifo_read/mem[11][1] ), .B(wdata_to_fifo[1]), .S0(n1210), 
        .Y(n279) );
  MX2 U1902 ( .A(\fifo_read/mem[11][2] ), .B(wdata_to_fifo[2]), .S0(n1210), 
        .Y(n278) );
  MX2 U1903 ( .A(\fifo_read/mem[11][3] ), .B(wdata_to_fifo[3]), .S0(n1210), 
        .Y(n277) );
  MX2 U1904 ( .A(\fifo_read/mem[11][4] ), .B(wdata_to_fifo[4]), .S0(n1210), 
        .Y(n276) );
  MX2 U1905 ( .A(\fifo_read/mem[11][5] ), .B(wdata_to_fifo[5]), .S0(n1210), 
        .Y(n275) );
  MX2 U1906 ( .A(\fifo_read/mem[11][6] ), .B(wdata_to_fifo[6]), .S0(n1210), 
        .Y(n274) );
  MX2 U1907 ( .A(\fifo_read/mem[11][7] ), .B(wdata_to_fifo[7]), .S0(n1210), 
        .Y(n273) );
  NOR2B U1908 ( .AN(n1428), .B(n1446), .Y(n1450) );
  MX2 U1909 ( .A(\fifo_read/mem[10][0] ), .B(n1316), .S0(n1212), .Y(n272) );
  MX2 U1910 ( .A(\fifo_read/mem[10][1] ), .B(n1314), .S0(n1212), .Y(n271) );
  MX2 U1911 ( .A(\fifo_read/mem[10][2] ), .B(n1328), .S0(n1212), .Y(n270) );
  MX2 U1912 ( .A(\fifo_read/mem[10][3] ), .B(n1326), .S0(n1212), .Y(n269) );
  MX2 U1913 ( .A(\fifo_read/mem[10][4] ), .B(n1324), .S0(n1212), .Y(n268) );
  MX2 U1914 ( .A(\fifo_read/mem[10][5] ), .B(n1322), .S0(n1212), .Y(n267) );
  MX2 U1915 ( .A(\fifo_read/mem[10][6] ), .B(n1336), .S0(n1212), .Y(n266) );
  MX2 U1916 ( .A(\fifo_read/mem[10][7] ), .B(n1334), .S0(n1212), .Y(n265) );
  NOR2B U1917 ( .AN(n1430), .B(n1446), .Y(n1451) );
  MX2 U1918 ( .A(\fifo_read/mem[9][0] ), .B(wdata_to_fifo[0]), .S0(n1190), .Y(
        n264) );
  MX2 U1919 ( .A(\fifo_read/mem[9][1] ), .B(wdata_to_fifo[1]), .S0(n1190), .Y(
        n263) );
  MX2 U1920 ( .A(\fifo_read/mem[9][2] ), .B(wdata_to_fifo[2]), .S0(n1190), .Y(
        n262) );
  MX2 U1921 ( .A(\fifo_read/mem[9][3] ), .B(wdata_to_fifo[3]), .S0(n1190), .Y(
        n261) );
  MX2 U1922 ( .A(\fifo_read/mem[9][4] ), .B(wdata_to_fifo[4]), .S0(n1190), .Y(
        n260) );
  MX2 U1923 ( .A(\fifo_read/mem[9][5] ), .B(wdata_to_fifo[5]), .S0(n1190), .Y(
        n259) );
  MX2 U1924 ( .A(\fifo_read/mem[9][6] ), .B(wdata_to_fifo[6]), .S0(n1190), .Y(
        n258) );
  MX2 U1925 ( .A(\fifo_read/mem[9][7] ), .B(wdata_to_fifo[7]), .S0(n1190), .Y(
        n257) );
  NOR2B U1926 ( .AN(n1432), .B(n1446), .Y(n1452) );
  MX2 U1927 ( .A(\fifo_read/mem[8][0] ), .B(n1316), .S0(n1192), .Y(n256) );
  MX2 U1928 ( .A(\fifo_read/mem[8][1] ), .B(n1314), .S0(n1192), .Y(n255) );
  MX2 U1929 ( .A(\fifo_read/mem[8][2] ), .B(n1328), .S0(n1192), .Y(n254) );
  MX2 U1930 ( .A(\fifo_read/mem[8][3] ), .B(n1326), .S0(n1192), .Y(n253) );
  MX2 U1931 ( .A(\fifo_read/mem[8][4] ), .B(n1324), .S0(n1192), .Y(n252) );
  MX2 U1932 ( .A(\fifo_read/mem[8][5] ), .B(n1322), .S0(n1192), .Y(n251) );
  MX2 U1933 ( .A(\fifo_read/mem[8][6] ), .B(n1336), .S0(n1192), .Y(n250) );
  MX2 U1934 ( .A(\fifo_read/mem[8][7] ), .B(n1334), .S0(n1192), .Y(n249) );
  NOR2B U1935 ( .AN(n1434), .B(n1446), .Y(n1453) );
  NAND3B U1936 ( .AN(\fifo_read/waddr[4] ), .B(n1435), .C(\fifo_read/waddr[3] ), .Y(n1446) );
  MX2 U1937 ( .A(\fifo_read/mem[7][0] ), .B(wdata_to_fifo[0]), .S0(n1194), .Y(
        n248) );
  MX2 U1938 ( .A(\fifo_read/mem[7][1] ), .B(wdata_to_fifo[1]), .S0(n1194), .Y(
        n247) );
  MX2 U1939 ( .A(\fifo_read/mem[7][2] ), .B(wdata_to_fifo[2]), .S0(n1194), .Y(
        n246) );
  MX2 U1940 ( .A(\fifo_read/mem[7][3] ), .B(wdata_to_fifo[3]), .S0(n1194), .Y(
        n245) );
  MX2 U1941 ( .A(\fifo_read/mem[7][4] ), .B(wdata_to_fifo[4]), .S0(n1194), .Y(
        n244) );
  MX2 U1942 ( .A(\fifo_read/mem[7][5] ), .B(wdata_to_fifo[5]), .S0(n1194), .Y(
        n243) );
  MX2 U1943 ( .A(\fifo_read/mem[7][6] ), .B(wdata_to_fifo[6]), .S0(n1194), .Y(
        n242) );
  MX2 U1944 ( .A(\fifo_read/mem[7][7] ), .B(wdata_to_fifo[7]), .S0(n1194), .Y(
        n241) );
  NOR2B U1945 ( .AN(n1419), .B(n1455), .Y(n1454) );
  NOR3B U1946 ( .AN(\fifo_read/waddr[2] ), .B(n1456), .C(n1457), .Y(n1419) );
  MX2 U1947 ( .A(\fifo_read/mem[6][0] ), .B(n1316), .S0(n1196), .Y(n240) );
  MX2 U1948 ( .A(\fifo_read/mem[6][1] ), .B(n1314), .S0(n1196), .Y(n239) );
  MX2 U1949 ( .A(\fifo_read/mem[6][2] ), .B(n1328), .S0(n1196), .Y(n238) );
  MX2 U1950 ( .A(\fifo_read/mem[6][3] ), .B(n1326), .S0(n1196), .Y(n237) );
  MX2 U1951 ( .A(\fifo_read/mem[6][4] ), .B(n1324), .S0(n1196), .Y(n236) );
  MX2 U1952 ( .A(\fifo_read/mem[6][5] ), .B(n1322), .S0(n1196), .Y(n235) );
  MX2 U1953 ( .A(\fifo_read/mem[6][6] ), .B(n1336), .S0(n1196), .Y(n234) );
  MX2 U1954 ( .A(\fifo_read/mem[6][7] ), .B(n1334), .S0(n1196), .Y(n233) );
  NOR2B U1955 ( .AN(n1422), .B(n1455), .Y(n1458) );
  NOR3B U1956 ( .AN(\fifo_read/waddr[2] ), .B(\fifo_read/waddr[0] ), .C(n1457), 
        .Y(n1422) );
  MX2 U1957 ( .A(\fifo_read/mem[5][0] ), .B(wdata_to_fifo[0]), .S0(n1198), .Y(
        n232) );
  MX2 U1958 ( .A(\fifo_read/mem[5][1] ), .B(wdata_to_fifo[1]), .S0(n1198), .Y(
        n231) );
  MX2 U1959 ( .A(\fifo_read/mem[5][2] ), .B(wdata_to_fifo[2]), .S0(n1198), .Y(
        n230) );
  MX2 U1960 ( .A(\fifo_read/mem[5][3] ), .B(wdata_to_fifo[3]), .S0(n1198), .Y(
        n229) );
  MX2 U1961 ( .A(\fifo_read/mem[5][4] ), .B(wdata_to_fifo[4]), .S0(n1198), .Y(
        n228) );
  MX2 U1962 ( .A(\fifo_read/mem[5][5] ), .B(wdata_to_fifo[5]), .S0(n1198), .Y(
        n227) );
  MX2 U1963 ( .A(\fifo_read/mem[5][6] ), .B(wdata_to_fifo[6]), .S0(n1198), .Y(
        n226) );
  MX2 U1964 ( .A(\fifo_read/mem[5][7] ), .B(wdata_to_fifo[7]), .S0(n1198), .Y(
        n225) );
  NOR2B U1965 ( .AN(n1424), .B(n1455), .Y(n1459) );
  NOR3B U1966 ( .AN(\fifo_read/waddr[2] ), .B(\fifo_read/waddr[1] ), .C(n1456), 
        .Y(n1424) );
  MX2 U1967 ( .A(\fifo_read/mem[4][0] ), .B(n1316), .S0(n1200), .Y(n224) );
  MX2 U1968 ( .A(\fifo_read/mem[4][1] ), .B(n1314), .S0(n1200), .Y(n223) );
  MX2 U1969 ( .A(\fifo_read/mem[4][2] ), .B(n1328), .S0(n1200), .Y(n222) );
  MX2 U1970 ( .A(\fifo_read/mem[4][3] ), .B(n1326), .S0(n1200), .Y(n221) );
  MX2 U1971 ( .A(\fifo_read/mem[4][4] ), .B(n1324), .S0(n1200), .Y(n220) );
  MX2 U1972 ( .A(\fifo_read/mem[4][5] ), .B(n1322), .S0(n1200), .Y(n219) );
  MX2 U1973 ( .A(\fifo_read/mem[4][6] ), .B(n1336), .S0(n1200), .Y(n218) );
  MX2 U1974 ( .A(\fifo_read/mem[4][7] ), .B(n1334), .S0(n1200), .Y(n217) );
  NOR2B U1975 ( .AN(n1426), .B(n1455), .Y(n1460) );
  NOR3B U1976 ( .AN(\fifo_read/waddr[2] ), .B(\fifo_read/waddr[0] ), .C(
        \fifo_read/waddr[1] ), .Y(n1426) );
  MX2 U1977 ( .A(\fifo_read/mem[3][0] ), .B(wdata_to_fifo[0]), .S0(n1202), .Y(
        n216) );
  MX2 U1978 ( .A(\fifo_read/mem[3][1] ), .B(wdata_to_fifo[1]), .S0(n1202), .Y(
        n215) );
  MX2 U1979 ( .A(\fifo_read/mem[3][2] ), .B(wdata_to_fifo[2]), .S0(n1202), .Y(
        n214) );
  MX2 U1980 ( .A(\fifo_read/mem[3][3] ), .B(wdata_to_fifo[3]), .S0(n1202), .Y(
        n213) );
  MX2 U1981 ( .A(\fifo_read/mem[3][4] ), .B(wdata_to_fifo[4]), .S0(n1202), .Y(
        n212) );
  MX2 U1982 ( .A(\fifo_read/mem[3][5] ), .B(wdata_to_fifo[5]), .S0(n1202), .Y(
        n211) );
  MX2 U1983 ( .A(\fifo_read/mem[3][6] ), .B(wdata_to_fifo[6]), .S0(n1202), .Y(
        n210) );
  MX2 U1984 ( .A(\fifo_read/mem[3][7] ), .B(wdata_to_fifo[7]), .S0(n1202), .Y(
        n209) );
  NOR2B U1985 ( .AN(n1428), .B(n1455), .Y(n1461) );
  NOR3 U1986 ( .A(\fifo_read/waddr[2] ), .B(n1456), .C(n1457), .Y(n1428) );
  MX2 U1987 ( .A(\fifo_read/mem[2][0] ), .B(n1316), .S0(n1204), .Y(n208) );
  MX2 U1988 ( .A(\fifo_read/mem[2][1] ), .B(n1314), .S0(n1204), .Y(n207) );
  MX2 U1989 ( .A(\fifo_read/mem[2][2] ), .B(n1328), .S0(n1204), .Y(n206) );
  MX2 U1990 ( .A(\fifo_read/mem[2][3] ), .B(n1326), .S0(n1204), .Y(n205) );
  MX2 U1991 ( .A(\fifo_read/mem[2][4] ), .B(n1324), .S0(n1204), .Y(n204) );
  MX2 U1992 ( .A(\fifo_read/mem[2][5] ), .B(n1322), .S0(n1204), .Y(n203) );
  MX2 U1993 ( .A(\fifo_read/mem[2][6] ), .B(n1336), .S0(n1204), .Y(n202) );
  MX2 U1994 ( .A(\fifo_read/mem[2][7] ), .B(n1334), .S0(n1204), .Y(n201) );
  NOR2B U1995 ( .AN(n1430), .B(n1455), .Y(n1462) );
  NOR3 U1996 ( .A(\fifo_read/waddr[2] ), .B(\fifo_read/waddr[0] ), .C(n1457), 
        .Y(n1430) );
  MX2 U1997 ( .A(\fifo_read/mem[1][0] ), .B(n1316), .S0(n1206), .Y(n200) );
  MX2 U1998 ( .A(\fifo_read/mem[1][1] ), .B(n1314), .S0(n1206), .Y(n199) );
  MX2 U1999 ( .A(\fifo_read/mem[1][2] ), .B(wdata_to_fifo[2]), .S0(n1206), .Y(
        n198) );
  MX2 U2000 ( .A(\fifo_read/mem[1][3] ), .B(wdata_to_fifo[3]), .S0(n1206), .Y(
        n197) );
  MX2 U2001 ( .A(\fifo_read/mem[1][4] ), .B(wdata_to_fifo[4]), .S0(n1206), .Y(
        n196) );
  MX2 U2002 ( .A(\fifo_read/mem[1][5] ), .B(wdata_to_fifo[5]), .S0(n1206), .Y(
        n195) );
  MX2 U2003 ( .A(\fifo_read/mem[1][6] ), .B(wdata_to_fifo[6]), .S0(n1206), .Y(
        n194) );
  MX2 U2004 ( .A(\fifo_read/mem[1][7] ), .B(n1334), .S0(n1206), .Y(n193) );
  NOR2B U2005 ( .AN(n1432), .B(n1455), .Y(n1463) );
  NOR2B U2006 ( .AN(n1464), .B(n1456), .Y(n1432) );
  MX2 U2007 ( .A(\fifo_read/mem[0][0] ), .B(n1316), .S0(n1208), .Y(n192) );
  MX2 U2008 ( .A(\fifo_read/mem[0][1] ), .B(n1314), .S0(n1208), .Y(n191) );
  MX2 U2009 ( .A(\fifo_read/mem[0][2] ), .B(n1328), .S0(n1208), .Y(n190) );
  MX2 U2010 ( .A(\fifo_read/mem[0][3] ), .B(n1326), .S0(n1208), .Y(n189) );
  MX2 U2011 ( .A(\fifo_read/mem[0][4] ), .B(n1324), .S0(n1208), .Y(n188) );
  MX2 U2012 ( .A(\fifo_read/mem[0][5] ), .B(n1322), .S0(n1208), .Y(n187) );
  MX2 U2013 ( .A(\fifo_read/mem[0][6] ), .B(n1336), .S0(n1208), .Y(n186) );
  MX2 U2014 ( .A(\fifo_read/mem[0][7] ), .B(n1334), .S0(n1208), .Y(n185) );
  NOR2B U2015 ( .AN(n1434), .B(n1455), .Y(n1465) );
  INV U2016 ( .A(n1466), .Y(n1455) );
  NOR3B U2017 ( .AN(n1435), .B(\fifo_read/waddr[4] ), .C(\fifo_read/waddr[3] ), 
        .Y(n1466) );
  NOR2B U2018 ( .AN(n1464), .B(\fifo_read/waddr[0] ), .Y(n1434) );
  NOR2 U2019 ( .A(\fifo_read/waddr[2] ), .B(\fifo_read/waddr[1] ), .Y(n1464)
         );
  NOR3B U2020 ( .AN(n1467), .B(n1468), .C(n1469), .Y(\fifo_write/wfull_next )
         );
  XNOR2 U2021 ( .A(\fifo_write/wbinnext[5] ), .B(\fifo_write/wq2_rgray [5]), 
        .Y(n1469) );
  XOR2 U2022 ( .A(\fifo_write/wgraynext[1] ), .B(\fifo_write/wq2_rgray [1]), 
        .Y(n1468) );
  XOR2 U2023 ( .A(\fifo_write/wbinnext[2] ), .B(\fifo_write/wbinnext[1] ), .Y(
        \fifo_write/wgraynext[1] ) );
  NOR4 U2024 ( .A(n1470), .B(n1471), .C(n1472), .D(n1473), .Y(n1467) );
  XNOR2 U2025 ( .A(\fifo_write/wgraynext[4] ), .B(\fifo_write/wq2_rgray [4]), 
        .Y(n1473) );
  XOR2 U2026 ( .A(\fifo_write/wbinnext[5] ), .B(\fifo_write/wbinnext[4] ), .Y(
        \fifo_write/wgraynext[4] ) );
  XOR2 U2027 ( .A(\fifo_write/wgraynext[2] ), .B(\fifo_write/wq2_rgray [2]), 
        .Y(n1472) );
  XOR2 U2028 ( .A(\fifo_write/wbinnext[3] ), .B(\fifo_write/wbinnext[2] ), .Y(
        \fifo_write/wgraynext[2] ) );
  XOR2 U2029 ( .A(\fifo_write/wgraynext[3] ), .B(\fifo_write/wq2_rgray [3]), 
        .Y(n1471) );
  XOR2 U2030 ( .A(\fifo_write/wbinnext[4] ), .B(\fifo_write/wbinnext[3] ), .Y(
        \fifo_write/wgraynext[3] ) );
  XOR2 U2031 ( .A(\fifo_write/wgraynext[0] ), .B(\fifo_write/wq2_rgray [0]), 
        .Y(n1470) );
  XOR2 U2032 ( .A(\fifo_write/wbinnext[1] ), .B(\fifo_write/wbinnext[0] ), .Y(
        \fifo_write/wgraynext[0] ) );
  XOR2 U2033 ( .A(\fifo_write/wgray [5]), .B(n1474), .Y(
        \fifo_write/wbinnext[5] ) );
  NOR2B U2034 ( .AN(\fifo_write/waddr[4] ), .B(n1475), .Y(n1474) );
  XNOR2 U2035 ( .A(\fifo_write/waddr[4] ), .B(n1475), .Y(
        \fifo_write/wbinnext[4] ) );
  NAND2 U2036 ( .A(\fifo_write/waddr[3] ), .B(n1476), .Y(n1475) );
  XOR2 U2037 ( .A(\fifo_write/waddr[3] ), .B(n1476), .Y(
        \fifo_write/wbinnext[3] ) );
  NOR2B U2038 ( .AN(n1477), .B(n1478), .Y(n1476) );
  INV U2039 ( .A(\fifo_write/waddr[2] ), .Y(n1478) );
  XOR2 U2040 ( .A(\fifo_write/waddr[2] ), .B(n1477), .Y(
        \fifo_write/wbinnext[2] ) );
  NOR2B U2041 ( .AN(n1479), .B(n1408), .Y(n1477) );
  INV U2042 ( .A(\fifo_write/waddr[1] ), .Y(n1408) );
  XOR2 U2043 ( .A(\fifo_write/waddr[1] ), .B(n1479), .Y(
        \fifo_write/wbinnext[1] ) );
  NOR2B U2044 ( .AN(n1386), .B(n1407), .Y(n1479) );
  INV U2045 ( .A(\fifo_write/waddr[0] ), .Y(n1407) );
  XOR2 U2046 ( .A(n1386), .B(\fifo_write/waddr[0] ), .Y(
        \fifo_write/wbinnext[0] ) );
  NOR2B U2047 ( .AN(i_wr), .B(fifo_1_w_full), .Y(n1386) );
  NOR4B U2048 ( .AN(n1480), .B(n1481), .C(n1482), .D(n1483), .Y(
        \fifo_write/rempty_next ) );
  XOR2 U2049 ( .A(\fifo_write/rgraynext[3] ), .B(\fifo_write/rq2_wgray [3]), 
        .Y(n1483) );
  XOR2 U2050 ( .A(\fifo_write/rbinnext[4] ), .B(\fifo_write/rbinnext[3] ), .Y(
        \fifo_write/rgraynext[3] ) );
  XOR2 U2051 ( .A(\fifo_write/rgraynext[1] ), .B(\fifo_write/rq2_wgray [1]), 
        .Y(n1482) );
  XOR2 U2052 ( .A(\fifo_write/rbinnext[2] ), .B(\fifo_write/rbinnext[1] ), .Y(
        \fifo_write/rgraynext[1] ) );
  XOR2 U2053 ( .A(\fifo_write/rbinnext[5] ), .B(\fifo_write/rq2_wgray [5]), 
        .Y(n1481) );
  NOR3 U2054 ( .A(n1484), .B(n1485), .C(n1486), .Y(n1480) );
  XOR2 U2055 ( .A(\fifo_write/rgraynext[2] ), .B(\fifo_write/rq2_wgray [2]), 
        .Y(n1486) );
  XOR2 U2056 ( .A(\fifo_write/rbinnext[3] ), .B(\fifo_write/rbinnext[2] ), .Y(
        \fifo_write/rgraynext[2] ) );
  XOR2 U2057 ( .A(\fifo_write/rgraynext[0] ), .B(\fifo_write/rq2_wgray [0]), 
        .Y(n1485) );
  XOR2 U2058 ( .A(\fifo_write/rbinnext[1] ), .B(\fifo_write/rbinnext[0] ), .Y(
        \fifo_write/rgraynext[0] ) );
  XOR2 U2059 ( .A(\fifo_write/rgraynext[4] ), .B(\fifo_write/rq2_wgray [4]), 
        .Y(n1484) );
  XOR2 U2060 ( .A(\fifo_write/rbinnext[5] ), .B(\fifo_write/rbinnext[4] ), .Y(
        \fifo_write/rgraynext[4] ) );
  XOR2 U2061 ( .A(\fifo_write/rgray [5]), .B(n1487), .Y(
        \fifo_write/rbinnext[5] ) );
  NOR2B U2062 ( .AN(n1188), .B(n1488), .Y(n1487) );
  XNOR2 U2063 ( .A(n1188), .B(n1488), .Y(\fifo_write/rbinnext[4] ) );
  NAND2 U2064 ( .A(n1489), .B(n1332), .Y(n1488) );
  XOR2 U2065 ( .A(n1489), .B(\fifo_write/rbin[3] ), .Y(
        \fifo_write/rbinnext[3] ) );
  NOR2B U2066 ( .AN(n1347), .B(n1490), .Y(n1489) );
  XNOR2 U2067 ( .A(n1348), .B(n1490), .Y(\fifo_write/rbinnext[2] ) );
  NAND2 U2068 ( .A(n1491), .B(n1341), .Y(n1490) );
  XOR2 U2069 ( .A(n1491), .B(n1183), .Y(\fifo_write/rbinnext[1] ) );
  NOR2B U2070 ( .AN(n1363), .B(n1492), .Y(n1491) );
  XNOR2 U2071 ( .A(n1360), .B(n1492), .Y(\fifo_write/rbinnext[0] ) );
  NAND2B U2072 ( .AN(rd_fifo_empty), .B(active), .Y(n1492) );
  NOR3B U2073 ( .AN(n1493), .B(n1494), .C(n1495), .Y(\fifo_read/wfull_next )
         );
  XNOR2 U2074 ( .A(\fifo_read/wbinnext[5] ), .B(\fifo_read/wq2_rgray [5]), .Y(
        n1495) );
  XOR2 U2075 ( .A(\fifo_read/wgraynext[1] ), .B(\fifo_read/wq2_rgray [1]), .Y(
        n1494) );
  XOR2 U2076 ( .A(\fifo_read/wbinnext[2] ), .B(\fifo_read/wbinnext[1] ), .Y(
        \fifo_read/wgraynext[1] ) );
  NOR4 U2077 ( .A(n1496), .B(n1497), .C(n1498), .D(n1499), .Y(n1493) );
  XNOR2 U2078 ( .A(\fifo_read/wgraynext[4] ), .B(\fifo_read/wq2_rgray [4]), 
        .Y(n1499) );
  XOR2 U2079 ( .A(\fifo_read/wbinnext[5] ), .B(\fifo_read/wbinnext[4] ), .Y(
        \fifo_read/wgraynext[4] ) );
  XOR2 U2080 ( .A(\fifo_read/wgraynext[2] ), .B(\fifo_read/wq2_rgray [2]), .Y(
        n1498) );
  XOR2 U2081 ( .A(\fifo_read/wbinnext[3] ), .B(\fifo_read/wbinnext[2] ), .Y(
        \fifo_read/wgraynext[2] ) );
  XOR2 U2082 ( .A(\fifo_read/wgraynext[3] ), .B(\fifo_read/wq2_rgray [3]), .Y(
        n1497) );
  XOR2 U2083 ( .A(\fifo_read/wbinnext[4] ), .B(\fifo_read/wbinnext[3] ), .Y(
        \fifo_read/wgraynext[3] ) );
  XOR2 U2084 ( .A(\fifo_read/wgraynext[0] ), .B(\fifo_read/wq2_rgray [0]), .Y(
        n1496) );
  XOR2 U2085 ( .A(\fifo_read/wbinnext[1] ), .B(\fifo_read/wbinnext[0] ), .Y(
        \fifo_read/wgraynext[0] ) );
  XOR2 U2086 ( .A(\fifo_read/wgray [5]), .B(n1500), .Y(\fifo_read/wbinnext[5] ) );
  NOR2B U2087 ( .AN(\fifo_read/waddr[4] ), .B(n1501), .Y(n1500) );
  XNOR2 U2088 ( .A(\fifo_read/waddr[4] ), .B(n1501), .Y(
        \fifo_read/wbinnext[4] ) );
  NAND2 U2089 ( .A(\fifo_read/waddr[3] ), .B(n1502), .Y(n1501) );
  XOR2 U2090 ( .A(\fifo_read/waddr[3] ), .B(n1502), .Y(\fifo_read/wbinnext[3] ) );
  NOR2B U2091 ( .AN(n1503), .B(n1504), .Y(n1502) );
  INV U2092 ( .A(\fifo_read/waddr[2] ), .Y(n1504) );
  XOR2 U2093 ( .A(\fifo_read/waddr[2] ), .B(n1503), .Y(\fifo_read/wbinnext[2] ) );
  NOR2B U2094 ( .AN(n1505), .B(n1457), .Y(n1503) );
  INV U2095 ( .A(\fifo_read/waddr[1] ), .Y(n1457) );
  XOR2 U2096 ( .A(\fifo_read/waddr[1] ), .B(n1505), .Y(\fifo_read/wbinnext[1] ) );
  NOR2B U2097 ( .AN(n1435), .B(n1456), .Y(n1505) );
  INV U2098 ( .A(\fifo_read/waddr[0] ), .Y(n1456) );
  XOR2 U2099 ( .A(n1435), .B(\fifo_read/waddr[0] ), .Y(\fifo_read/wbinnext[0] ) );
  NOR2B U2100 ( .AN(active), .B(o_wfull), .Y(n1435) );
  NOR4B U2101 ( .AN(n1506), .B(n1507), .C(n1508), .D(n1509), .Y(
        \fifo_read/rempty_next ) );
  XOR2 U2102 ( .A(\fifo_read/rgraynext[3] ), .B(\fifo_read/rq2_wgray [3]), .Y(
        n1509) );
  XOR2 U2103 ( .A(\fifo_read/rbinnext[4] ), .B(\fifo_read/rbinnext[3] ), .Y(
        \fifo_read/rgraynext[3] ) );
  XOR2 U2104 ( .A(\fifo_read/rgraynext[1] ), .B(\fifo_read/rq2_wgray [1]), .Y(
        n1508) );
  XOR2 U2105 ( .A(\fifo_read/rbinnext[2] ), .B(\fifo_read/rbinnext[1] ), .Y(
        \fifo_read/rgraynext[1] ) );
  XOR2 U2106 ( .A(\fifo_read/rbinnext[5] ), .B(\fifo_read/rq2_wgray [5]), .Y(
        n1507) );
  NOR3 U2107 ( .A(n1510), .B(n1511), .C(n1512), .Y(n1506) );
  XOR2 U2108 ( .A(\fifo_read/rgraynext[2] ), .B(\fifo_read/rq2_wgray [2]), .Y(
        n1512) );
  XOR2 U2109 ( .A(\fifo_read/rbinnext[3] ), .B(\fifo_read/rbinnext[2] ), .Y(
        \fifo_read/rgraynext[2] ) );
  XOR2 U2110 ( .A(\fifo_read/rgraynext[0] ), .B(\fifo_read/rq2_wgray [0]), .Y(
        n1511) );
  XOR2 U2111 ( .A(\fifo_read/rbinnext[1] ), .B(\fifo_read/rbinnext[0] ), .Y(
        \fifo_read/rgraynext[0] ) );
  XOR2 U2112 ( .A(\fifo_read/rgraynext[4] ), .B(\fifo_read/rq2_wgray [4]), .Y(
        n1510) );
  XOR2 U2113 ( .A(\fifo_read/rbinnext[5] ), .B(\fifo_read/rbinnext[4] ), .Y(
        \fifo_read/rgraynext[4] ) );
  XOR2 U2114 ( .A(\fifo_read/rgray [5]), .B(n1513), .Y(\fifo_read/rbinnext[5] ) );
  NOR2B U2115 ( .AN(n1186), .B(n1514), .Y(n1513) );
  XNOR2 U2116 ( .A(n1186), .B(n1514), .Y(\fifo_read/rbinnext[4] ) );
  NAND2 U2117 ( .A(n1515), .B(n1330), .Y(n1514) );
  XOR2 U2118 ( .A(n1515), .B(\fifo_read/rbin[3] ), .Y(\fifo_read/rbinnext[3] )
         );
  NOR2B U2119 ( .AN(n1344), .B(n1516), .Y(n1515) );
  XNOR2 U2120 ( .A(n1345), .B(n1516), .Y(\fifo_read/rbinnext[2] ) );
  NAND2 U2121 ( .A(n1517), .B(n1338), .Y(n1516) );
  XOR2 U2122 ( .A(n1517), .B(n1181), .Y(\fifo_read/rbinnext[1] ) );
  NOR2B U2123 ( .AN(n1353), .B(n1518), .Y(n1517) );
  XNOR2 U2124 ( .A(n1350), .B(n1518), .Y(\fifo_read/rbinnext[0] ) );
  NAND2B U2125 ( .AN(o_rempty), .B(i_rd), .Y(n1518) );
  NOR2 U2126 ( .A(rd_fifo_empty), .B(rst), .Y(N2) );
endmodule
